`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:48:10 12/03/2013 
// Design Name: 
// Module Name:    des_translate 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module des_translate(clk, rst, flag, ready, datain, key, dataout);
input clk;
  input rst;
  input flag;
  output ready;
  input [64 : 1] datain;
  input [64 : 1] key;
  output [64 : 1] dataout;
  wire clk_BUFGP;
  wire rst_IBUF;
  wire flag_IBUF;
  wire N5008;
  wire ready_OBUF;
  wire \MUX_BLOCK_roundsel<1>_mmx_out55 ;
  wire \MUX_BLOCK_roundsel<2>_mmx_out27 ;
  wire CHOICE1134;
  wire \c1/u4/Mrom_dout_N6 ;
  wire \c1/u5/Mrom_dout_N6 ;
  wire _n0000;
  wire _n0001;
  wire state_FFd4;
  wire state_FFd2;
  wire state_FFd1;
  wire state_FFd7;
  wire N5009;
  wire state_FFd6;
  wire state_FFd5;
  wire state_FFd8;
  wire state_FFd3;
  wire N5897;
  wire \c1/u3/Mrom_dout_inst_lut4_78 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out68 ;
  wire \c1/u3/Mrom_dout_inst_lut4_76 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out70 ;
  wire \c1/u3/Mrom_dout_N9 ;
  wire _n0030;
  wire _n0025;
  wire \MUX_BLOCK_roundsel<1>_mmx_out48 ;
  wire \c1/u5/Mrom_dout_N1 ;
  wire \c1/u5/Mrom_dout_inst_lut4_43 ;
  wire \c1/u5/Mrom_dout_inst_lut4_37 ;
  wire \c1/u5/Mrom_dout_N9 ;
  wire _n0029;
  wire \key1[4] ;
  wire \c1/u5/Mrom_dout_inst_lut4_46 ;
  wire \key1[5] ;
  wire \c1/u5/Mrom_dout_inst_lut4_44 ;
  wire \key1[6] ;
  wire N5011;
  wire \key1[7] ;
  wire \key1[2] ;
  wire \key1[8] ;
  wire \key1[3] ;
  wire \key1[64] ;
  wire \key1[14] ;
  wire \state_FFd6-In ;
  wire \c1/u4/Mrom_dout_N1 ;
  wire \key1[15] ;
  wire \key1[10] ;
  wire \c1/u4/Mrom_dout_inst_lut4_53 ;
  wire \key1[16] ;
  wire \key1[11] ;
  wire \c1/u4/Mrom_dout_inst_lut4_55 ;
  wire \state_FFd3-In ;
  wire \key1[12] ;
  wire N1;
  wire \key1[18] ;
  wire \key1[13] ;
  wire CHOICE1038;
  wire \key1[24] ;
  wire \key1[19] ;
  wire CHOICE900;
  wire \MUX_BLOCK_roundsel<1>_mmx_out6 ;
  wire \key1[20] ;
  wire \c1/u3/Mrom_dout_inst_lut4_75 ;
  wire \key1[26] ;
  wire \key1[21] ;
  wire \key1[27] ;
  wire \key1[22] ;
  wire \key1[28] ;
  wire \key1[23] ;
  wire \key1[34] ;
  wire \key1[29] ;
  wire \key1[35] ;
  wire \key1[30] ;
  wire \key1[36] ;
  wire \key1[31] ;
  wire \key1[37] ;
  wire \key1[32] ;
  wire \key1[38] ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out7 ;
  wire \key1[44] ;
  wire \key1[39] ;
  wire \key1[45] ;
  wire \key1[40] ;
  wire \key1[46] ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out69 ;
  wire \key1[47] ;
  wire \key1[42] ;
  wire \key1[48] ;
  wire \key1[43] ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out10 ;
  wire \key1[54] ;
  wire \state_FFd5-In ;
  wire \key1[55] ;
  wire \key1[50] ;
  wire \key1[56] ;
  wire \key1[51] ;
  wire \c1/u3/Mrom_dout_inst_lut4_65 ;
  wire \key1[52] ;
  wire \key1[58] ;
  wire \key1[53] ;
  wire \key1[59] ;
  wire N5010;
  wire \key1[60] ;
  wire \key1[61] ;
  wire \key1[62] ;
  wire \key1[63] ;
  wire \c1/u5/Mrom_dout_inst_lut4_35 ;
  wire dataout_64;
  wire dataout_63;
  wire dataout_62;
  wire dataout_61;
  wire dataout_60;
  wire dataout_59;
  wire dataout_58;
  wire dataout_57;
  wire dataout_56;
  wire dataout_55;
  wire dataout_54;
  wire dataout_53;
  wire dataout_52;
  wire dataout_51;
  wire dataout_50;
  wire dataout_49;
  wire dataout_48;
  wire dataout_47;
  wire dataout_46;
  wire dataout_45;
  wire dataout_44;
  wire dataout_43;
  wire dataout_42;
  wire dataout_41;
  wire dataout_40;
  wire dataout_39;
  wire dataout_38;
  wire dataout_37;
  wire dataout_36;
  wire dataout_35;
  wire dataout_34;
  wire dataout_33;
  wire dataout_32;
  wire dataout_31;
  wire dataout_30;
  wire dataout_29;
  wire dataout_28;
  wire dataout_27;
  wire dataout_26;
  wire dataout_25;
  wire dataout_24;
  wire dataout_23;
  wire dataout_22;
  wire dataout_21;
  wire dataout_20;
  wire dataout_19;
  wire dataout_18;
  wire dataout_17;
  wire dataout_16;
  wire dataout_15;
  wire dataout_14;
  wire dataout_13;
  wire dataout_12;
  wire dataout_11;
  wire dataout_10;
  wire dataout_9;
  wire dataout_8;
  wire dataout_7;
  wire dataout_6;
  wire dataout_5;
  wire dataout_4;
  wire dataout_3;
  wire dataout_2;
  wire dataout_1;
  wire datain_64_IBUF;
  wire datain_63_IBUF;
  wire datain_62_IBUF;
  wire datain_61_IBUF;
  wire datain_60_IBUF;
  wire datain_59_IBUF;
  wire datain_58_IBUF;
  wire datain_57_IBUF;
  wire datain_56_IBUF;
  wire datain_55_IBUF;
  wire datain_54_IBUF;
  wire datain_53_IBUF;
  wire datain_52_IBUF;
  wire datain_51_IBUF;
  wire datain_50_IBUF;
  wire datain_49_IBUF;
  wire datain_48_IBUF;
  wire datain_47_IBUF;
  wire datain_46_IBUF;
  wire datain_45_IBUF;
  wire datain_44_IBUF;
  wire datain_43_IBUF;
  wire datain_42_IBUF;
  wire datain_41_IBUF;
  wire datain_40_IBUF;
  wire datain_39_IBUF;
  wire datain_38_IBUF;
  wire datain_37_IBUF;
  wire datain_36_IBUF;
  wire datain_35_IBUF;
  wire datain_34_IBUF;
  wire datain_33_IBUF;
  wire datain_32_IBUF;
  wire datain_31_IBUF;
  wire datain_30_IBUF;
  wire datain_29_IBUF;
  wire datain_28_IBUF;
  wire datain_27_IBUF;
  wire datain_26_IBUF;
  wire datain_25_IBUF;
  wire datain_24_IBUF;
  wire datain_23_IBUF;
  wire datain_22_IBUF;
  wire datain_21_IBUF;
  wire datain_20_IBUF;
  wire datain_19_IBUF;
  wire datain_18_IBUF;
  wire datain_17_IBUF;
  wire datain_16_IBUF;
  wire datain_15_IBUF;
  wire datain_14_IBUF;
  wire datain_13_IBUF;
  wire datain_12_IBUF;
  wire datain_11_IBUF;
  wire datain_10_IBUF;
  wire datain_9_IBUF;
  wire datain_8_IBUF;
  wire datain_7_IBUF;
  wire datain_6_IBUF;
  wire datain_5_IBUF;
  wire datain_4_IBUF;
  wire datain_3_IBUF;
  wire datain_2_IBUF;
  wire datain_1_IBUF;
  wire key_64_IBUF;
  wire key_63_IBUF;
  wire key_62_IBUF;
  wire key_61_IBUF;
  wire key_60_IBUF;
  wire key_59_IBUF;
  wire key_58_IBUF;
  wire \c1/u3/Mrom_dout_inst_lut4_67 ;
  wire key_56_IBUF;
  wire key_55_IBUF;
  wire key_54_IBUF;
  wire key_53_IBUF;
  wire key_52_IBUF;
  wire key_51_IBUF;
  wire key_50_IBUF;
  wire key_48_IBUF;
  wire key_47_IBUF;
  wire key_46_IBUF;
  wire key_45_IBUF;
  wire key_44_IBUF;
  wire key_43_IBUF;
  wire key_42_IBUF;
  wire key_40_IBUF;
  wire key_39_IBUF;
  wire key_38_IBUF;
  wire key_37_IBUF;
  wire key_36_IBUF;
  wire key_35_IBUF;
  wire key_34_IBUF;
  wire key_32_IBUF;
  wire key_31_IBUF;
  wire key_30_IBUF;
  wire key_29_IBUF;
  wire key_28_IBUF;
  wire key_27_IBUF;
  wire key_26_IBUF;
  wire key_24_IBUF;
  wire key_23_IBUF;
  wire key_22_IBUF;
  wire key_21_IBUF;
  wire key_20_IBUF;
  wire key_19_IBUF;
  wire key_18_IBUF;
  wire key_16_IBUF;
  wire key_15_IBUF;
  wire key_14_IBUF;
  wire key_13_IBUF;
  wire key_12_IBUF;
  wire key_11_IBUF;
  wire key_10_IBUF;
  wire key_8_IBUF;
  wire key_7_IBUF;
  wire key_6_IBUF;
  wire key_5_IBUF;
  wire key_4_IBUF;
  wire key_3_IBUF;
  wire key_2_IBUF;
  wire N5087;
  wire N5085;
  wire N5089;
  wire N5091;
  wire N5153;
  wire \key2[7] ;
  wire N5093;
  wire N5059;
  wire N5061;
  wire N5171;
  wire N5115;
  wire N5063;
  wire N5095;
  wire N5097;
  wire N5179;
  wire \key2[19] ;
  wire N5065;
  wire N5099;
  wire N5067;
  wire N5069;
  wire N5123;
  wire N5117;
  wire N5101;
  wire N5103;
  wire N5071;
  wire N5155;
  wire \key2[31] ;
  wire N5073;
  wire N5075;
  wire N5105;
  wire N5157;
  wire N5119;
  wire N5077;
  wire N5107;
  wire N5109;
  wire N5079;
  wire N5125;
  wire N5121;
  wire N5081;
  wire N5111;
  wire N5113;
  wire N5083;
  wire N5159;
  wire \c1/u5/Mrom_dout_inst_lut4_33 ;
  wire \c1/u5/Mrom_dout_inst_lut4_39 ;
  wire \c1/u5/Mrom_dout_inst_lut4_41 ;
  wire CHOICE1268;
  wire \c1/u4/Mrom_dout_inst_lut4_60 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out8 ;
  wire \c1/u5/Mrom_dout_N4 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out67 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out9 ;
  wire \c1/u4/Mrom_dout_inst_lut4_62 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out46 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out45 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out50 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out49 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out95 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out94 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out63 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out93 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out92 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out91 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out62 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out90 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out44 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out43 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out42 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out41 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out40 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out39 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out38 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out37 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out36 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out35 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out34 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out33 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out32 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out51 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out47 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out31 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out30 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out29 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out28 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out27 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out1 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out26 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out25 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out2 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out24 ;
  wire N01;
  wire \MUX_BLOCK_roundsel<1>_mmx_out23 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out3 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out22 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out21 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out5 ;
  wire \MUX_BLOCK_roundsel<2>_mmx_out11 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out4 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out66 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out20 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out65 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out19 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out18 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out17 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out16 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out15 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out14 ;
  wire \MUX_BLOCK_roundsel<2>_mmx_out7 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out13 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out64 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out12 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out11 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out89 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out88 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out87 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out86 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out85 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out61 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out84 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out83 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out82 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out81 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out80 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out79 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out54 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out78 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out60 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out59 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out58 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out77 ;
  wire \MUX_BLOCK_roundsel<2>_mmx_out33 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out53 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out76 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out75 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out74 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out73 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out57 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out56 ;
  wire \MUX_BLOCK_roundsel<2>_mmx_out24 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out72 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out52 ;
  wire \MUX_BLOCK_roundsel<1>_mmx_out71 ;
  wire \c1/u5/Mrom_dout_N10 ;
  wire \c1/u5/Mrom_dout_inst_lut4_42 ;
  wire \c1/X[1] ;
  wire \c1/u3/Mrom_dout_inst_lut4_71 ;
  wire \c1/u5/Mrom_dout_inst_lut4_47 ;
  wire N5175;
  wire \c1/u3/Mrom_dout_inst_lut4_72 ;
  wire \c1/u3/Mrom_dout_inst_lut4_73 ;
  wire \c1/u2/Mrom_dout_inst_lut4_90 ;
  wire \c1/u2/Mrom_dout_inst_lut4_91 ;
  wire \c1/X[8] ;
  wire \c1/X[6] ;
  wire \c1/X[4] ;
  wire \c1/X[2] ;
  wire \c1/X[48] ;
  wire \c1/X[10] ;
  wire \c1/X[37] ;
  wire \c1/u2/Mrom_dout_inst_lut4_95 ;
  wire \c1/X[11] ;
  wire \c1/u5/Mrom_dout_N0 ;
  wire \c1/u3/Mrom_dout_N10 ;
  wire \c1/X[18] ;
  wire \c1/u4/Mrom_dout_inst_lut4_61 ;
  wire \c1/X[20] ;
  wire \c1/u5/Mrom_dout_N7 ;
  wire \c1/X[22] ;
  wire CHOICE1954;
  wire \c1/X[24] ;
  wire \c1/u3/Mrom_dout_inst_lut4_66 ;
  wire \c1/u5/Mrom_dout_inst_lut4_38 ;
  wire \c1/X[17] ;
  wire \c1/X[38] ;
  wire \c1/X[28] ;
  wire \c1/X[40] ;
  wire \c1/X[30] ;
  wire \c1/X[42] ;
  wire \c1/X[32] ;
  wire \c1/u2/Mrom_dout_inst_lut4_94 ;
  wire \c1/X[44] ;
  wire \c1/X[34] ;
  wire \c1/X[25] ;
  wire \c1/X[27] ;
  wire \c1/X[15] ;
  wire \c1/X[12] ;
  wire \c1/u3/Mrom_dout_inst_lut4_74 ;
  wire \c1/X[47] ;
  wire \c1/u5/Mrom_dout_inst_lut4_45 ;
  wire \c1/u4/Mrom_dout_inst_lut4_52 ;
  wire \c1/u4/Mrom_dout_N7 ;
  wire \c1/u5/Mrom_dout_N3 ;
  wire N5151;
  wire \c1/u3/Mrom_dout_inst_lut4_64 ;
  wire \c1/u5/Mrom_dout_inst_lut4_34 ;
  wire \c1/u5/Mrom_dout_inst_lut4_36 ;
  wire CHOICE1162;
  wire \c1/u5/Mrom_dout_inst_lut4_40 ;
  wire \c1/u5/Mrom_dout_inst_lut4_32 ;
  wire \c1/u4/Mrom_dout_N0 ;
  wire \c1/u3/Mrom_dout_inst_lut4_69 ;
  wire \c1/u4/Mrom_dout_inst_lut4_63 ;
  wire CHOICE1955;
  wire \c1/X[35] ;
  wire \c1/X[45] ;
  wire \c1/X[14] ;
  wire \c1/X[46] ;
  wire \c1/X[43] ;
  wire \c1/X[41] ;
  wire \c1/X[39] ;
  wire \c1/X[36] ;
  wire \c1/X[33] ;
  wire \c1/X[29] ;
  wire \c1/X[26] ;
  wire \c1/X[23] ;
  wire \c1/X[21] ;
  wire \c1/X[19] ;
  wire \c1/X[16] ;
  wire CHOICE1405;
  wire CHOICE1340;
  wire \c1/u4/Mrom_dout_inst_lut4_54 ;
  wire \c1/X[13] ;
  wire \c1/u2/Mrom_dout_inst_lut4_93 ;
  wire \c1/u2/Mrom_dout_inst_lut4_92 ;
  wire \c1/X[3] ;
  wire \c1/X[5] ;
  wire \c1/X[9] ;
  wire \c1/u6/Mrom_dout_inst_lut4_25 ;
  wire \c1/u6/Mrom_dout_inst_lut4_24 ;
  wire \c1/u6/Mrom_dout_N4 ;
  wire \c1/u6/Mrom_dout_N3 ;
  wire N5448;
  wire CHOICE1029;
  wire \c1/u6/Mrom_dout_inst_lut4_19 ;
  wire \c1/u6/Mrom_dout_inst_lut4_18 ;
  wire \c1/u6/Mrom_dout_inst_lut4_17 ;
  wire \c1/u6/Mrom_dout_inst_lut4_16 ;
  wire CHOICE1615;
  wire \c1/u6/Mrom_dout_inst_lut4_29 ;
  wire \c1/u6/Mrom_dout_inst_lut4_30 ;
  wire \c1/u6/Mrom_dout_inst_lut4_31 ;
  wire CHOICE1897;
  wire \c1/u6/Mrom_dout_inst_lut4_27 ;
  wire \c1/u6/Mrom_dout_inst_lut4_26 ;
  wire \c1/u7/Mrom_dout_inst_lut4_11 ;
  wire \c1/u7/Mrom_dout_inst_lut4_10 ;
  wire N5490;
  wire CHOICE1267;
  wire \c1/u7/Mrom_dout_inst_lut4_7 ;
  wire \c1/u7/Mrom_dout_inst_lut4_6 ;
  wire \c1/u1/Mrom_dout_inst_lut4_121 ;
  wire \c1/u1/Mrom_dout_inst_lut4_120 ;
  wire \c1/u1/Mrom_dout_N4 ;
  wire \c1/u1/Mrom_dout_N3 ;
  wire \c1/u1/Mrom_dout_inst_lut4_119 ;
  wire \c1/u1/Mrom_dout_inst_lut4_118 ;
  wire \c1/u1/Mrom_dout_inst_lut4_117 ;
  wire \c1/u1/Mrom_dout_inst_lut4_116 ;
  wire \c1/u1/Mrom_dout_N1 ;
  wire \c1/u1/Mrom_dout_N0 ;
  wire \c1/u1/Mrom_dout_inst_lut4_115 ;
  wire \c1/u1/Mrom_dout_inst_lut4_114 ;
  wire \c1/u1/Mrom_dout_inst_lut4_113 ;
  wire \c1/u1/Mrom_dout_inst_lut4_112 ;
  wire \c1/u1/Mrom_dout_N6 ;
  wire \c1/u1/Mrom_dout_N7 ;
  wire N5187;
  wire N5186;
  wire N5184;
  wire N5183;
  wire \c1/u1/Mrom_dout_N9 ;
  wire \c1/u1/Mrom_dout_N10 ;
  wire \c1/u1/Mrom_dout_inst_lut4_123 ;
  wire \c1/u1/Mrom_dout_inst_lut4_122 ;
  wire \c1/u0/Mrom_dout_inst_lut4_105 ;
  wire \c1/u0/Mrom_dout_inst_lut4_104 ;
  wire CHOICE1833;
  wire CHOICE1332;
  wire \c1/u0/Mrom_dout_inst_lut4_103 ;
  wire \c1/u0/Mrom_dout_inst_lut4_102 ;
  wire \c1/u0/Mrom_dout_inst_lut4_101 ;
  wire \c1/u0/Mrom_dout_inst_lut4_100 ;
  wire N5035;
  wire CHOICE1320;
  wire \c1/u0/Mrom_dout_inst_lut4_99 ;
  wire \c1/u0/Mrom_dout_inst_lut4_98 ;
  wire \c1/u0/Mrom_dout_inst_lut4_97 ;
  wire \c1/u0/Mrom_dout_inst_lut4_96 ;
  wire CHOICE1206;
  wire \c1/u0/Mrom_dout_inst_lut4_108 ;
  wire \c1/u0/Mrom_dout_inst_lut4_109 ;
  wire \c1/u0/Mrom_dout_inst_lut4_110 ;
  wire \c1/u0/Mrom_dout_inst_lut4_111 ;
  wire N5047;
  wire CHOICE1553;
  wire \c1/u0/Mrom_dout_inst_lut4_107 ;
  wire \c1/u0/Mrom_dout_inst_lut4_106 ;
  wire \c1/u2/Mrom_dout_inst_lut4_89 ;
  wire \c1/u2/Mrom_dout_inst_lut4_88 ;
  wire N5430;
  wire \c1/u2/Mrom_dout_inst_lut4_87 ;
  wire \c1/u2/Mrom_dout_inst_lut4_86 ;
  wire \c1/u2/Mrom_dout_inst_lut4_85 ;
  wire \c1/u2/Mrom_dout_inst_lut4_84 ;
  wire N5181;
  wire \c1/u2/Mrom_dout_inst_lut4_83 ;
  wire \c1/u2/Mrom_dout_inst_lut4_82 ;
  wire \c1/u2/Mrom_dout_inst_lut4_81 ;
  wire \c1/u2/Mrom_dout_inst_lut4_80 ;
  wire \c1/u7/Mrom_dout_inst_lut4_4 ;
  wire \c1/u7/Mrom_dout_inst_lut4_5 ;
  wire N5482;
  wire \c1/u7/Mrom_dout_inst_lut4_15 ;
  wire \c1/u7/Mrom_dout_inst_lut4_14 ;
  wire \c1/u7/Mrom_dout_inst_lut4_13 ;
  wire \c1/u7/Mrom_dout_inst_lut4_12 ;
  wire CHOICE1011;
  wire \c1/u7/Mrom_dout_inst_lut4_0 ;
  wire \c1/u7/Mrom_dout_inst_lut4_1 ;
  wire \c1/u7/Mrom_dout_inst_lut4_2 ;
  wire \c1/u7/Mrom_dout_inst_lut4_3 ;
  wire CHOICE1918;
  wire N234;
  wire CHOICE1652;
  wire CHOICE13;
  wire CHOICE1936;
  wire CHOICE2;
  wire CHOICE740;
  wire CHOICE195;
  wire CHOICE503;
  wire CHOICE734;
  wire CHOICE23;
  wire CHOICE19;
  wire N5484;
  wire CHOICE1928;
  wire CHOICE136;
  wire CHOICE311;
  wire CHOICE831;
  wire CHOICE21;
  wire CHOICE678;
  wire CHOICE497;
  wire CHOICE149;
  wire CHOICE32;
  wire CHOICE531;
  wire CHOICE936;
  wire CHOICE824;
  wire CHOICE28;
  wire N5446;
  wire N5033;
  wire CHOICE423;
  wire CHOICE145;
  wire CHOICE463;
  wire CHOICE30;
  wire CHOICE140;
  wire CHOICE822;
  wire CHOICE138;
  wire CHOICE964;
  wire CHOICE41;
  wire CHOICE819;
  wire CHOICE147;
  wire CHOICE611;
  wire CHOICE1104;
  wire CHOICE37;
  wire CHOICE1645;
  wire N5444;
  wire CHOICE475;
  wire CHOICE339;
  wire CHOICE39;
  wire CHOICE731;
  wire CHOICE733;
  wire CHOICE50;
  wire N5476;
  wire CHOICE1086;
  wire CHOICE1823;
  wire CHOICE46;
  wire CHOICE510;
  wire N5452;
  wire CHOICE156;
  wire CHOICE675;
  wire CHOICE158;
  wire CHOICE48;
  wire CHOICE812;
  wire N5456;
  wire CHOICE367;
  wire CHOICE59;
  wire N5488;
  wire CHOICE283;
  wire N5141;
  wire CHOICE1234;
  wire CHOICE55;
  wire CHOICE1046;
  wire N5466;
  wire CHOICE722;
  wire CHOICE57;
  wire CHOICE154;
  wire CHOICE803;
  wire CHOICE68;
  wire CHOICE1927;
  wire CHOICE230;
  wire N5129;
  wire N5133;
  wire CHOICE64;
  wire CHOICE660;
  wire N5195;
  wire CHOICE794;
  wire CHOICE66;
  wire N5474;
  wire N5499;
  wire N5440;
  wire CHOICE785;
  wire CHOICE77;
  wire N5454;
  wire CHOICE713;
  wire CHOICE73;
  wire CHOICE616;
  wire CHOICE651;
  wire CHOICE788;
  wire CHOICE75;
  wire CHOICE399;
  wire CHOICE633;
  wire CHOICE787;
  wire CHOICE86;
  wire CHOICE1047;
  wire N5464;
  wire N5460;
  wire CHOICE82;
  wire CHOICE259;
  wire N5495;
  wire N5472;
  wire CHOICE84;
  wire CHOICE1789;
  wire N5199;
  wire CHOICE626;
  wire N5442;
  wire CHOICE95;
  wire CHOICE642;
  wire CHOICE1913;
  wire CHOICE1122;
  wire CHOICE91;
  wire N5500;
  wire CHOICE776;
  wire CHOICE391;
  wire CHOICE93;
  wire CHOICE595;
  wire CHOICE104;
  wire CHOICE686;
  wire CHOICE767;
  wire CHOICE455;
  wire CHOICE100;
  wire CHOICE704;
  wire CHOICE585;
  wire CHOICE102;
  wire CHOICE695;
  wire CHOICE113;
  wire N5450;
  wire CHOICE758;
  wire CHOICE109;
  wire CHOICE431;
  wire N5470;
  wire CHOICE521;
  wire CHOICE579;
  wire CHOICE111;
  wire CHOICE1849;
  wire CHOICE491;
  wire CHOICE122;
  wire CHOICE1262;
  wire CHOICE1106;
  wire CHOICE751;
  wire CHOICE680;
  wire CHOICE118;
  wire N5462;
  wire CHOICE669;
  wire N5458;
  wire CHOICE199;
  wire CHOICE120;
  wire CHOICE624;
  wire CHOICE749;
  wire CHOICE752;
  wire CHOICE131;
  wire N5428;
  wire CHOICE1437;
  wire N5468;
  wire CHOICE127;
  wire CHOICE547;
  wire CHOICE571;
  wire CHOICE129;
  wire CHOICE2017;
  wire N5478;
  wire N5432;
  wire CHOICE1817;
  wire CHOICE840;
  wire CHOICE1178;
  wire N5139;
  wire CHOICE1887;
  wire CHOICE1310;
  wire CHOICE867;
  wire CHOICE2008;
  wire CHOICE1190;
  wire CHOICE1277;
  wire N5135;
  wire N5017;
  wire CHOICE1705;
  wire CHOICE1855;
  wire CHOICE849;
  wire CHOICE1074;
  wire CHOICE970;
  wire CHOICE2009;
  wire CHOICE851;
  wire N5173;
  wire CHOICE1639;
  wire CHOICE1733;
  wire N5438;
  wire N5177;
  wire CHOICE1377;
  wire CHOICE1609;
  wire N5039;
  wire CHOICE1411;
  wire CHOICE1304;
  wire N5436;
  wire CHOICE1621;
  wire CHOICE1663;
  wire CHOICE1999;
  wire CHOICE1577;
  wire CHOICE1761;
  wire CHOICE1990;
  wire CHOICE1545;
  wire CHOICE1150;
  wire CHOICE1056;
  wire N5486;
  wire CHOICE1981;
  wire CHOICE1982;
  wire CHOICE1521;
  wire CHOICE873;
  wire CHOICE1465;
  wire CHOICE1080;
  wire N5131;
  wire CHOICE1276;
  wire CHOICE1020;
  wire N5169;
  wire N5193;
  wire CHOICE1002;
  wire CHOICE1945;
  wire CHOICE1964;
  wire N5045;
  wire CHOICE1881;
  wire CHOICE1093;
  wire N5019;
  wire CHOICE1973;
  wire N5021;
  wire CHOICE1946;
  wire CHOICE1972;
  wire CHOICE1676;
  wire CHOICE1058;
  wire CHOICE1669;
  wire CHOICE1345;
  wire N5434;
  wire CHOICE908;
  wire N5480;
  wire CHOICE1865;
  wire CHOICE996;
  wire CHOICE1937;
  wire CHOICE1963;
  wire CHOICE1585;
  wire CHOICE1493;
  wire CHOICE1421;
  wire CHOICE1628;
  wire CHOICE980;
  wire N5137;
  wire roundsel_11;
  wire roundsel_3_1;
  wire roundsel_2_1;
  wire roundsel_4_1;
  wire Ker039;
  wire roundsel_1_1;
  wire roundsel_32;
  wire roundsel_22;
  wire roundsel_12;
  wire roundsel_4_2;
  wire roundsel_1_11;
  wire roundsel_1_3;
  wire roundsel_1_6;
  wire roundsel_23;
  wire roundsel_33;
  wire roundsel_43;
  wire roundsel_2_4;
  wire roundsel_3_2;
  wire roundsel_1_2;
  wire roundsel_1_4;
  wire roundsel_1_5;
  wire roundsel_1_10;
  wire roundsel_3_3;
  wire roundsel_4_3;
  wire roundsel_24;
  wire roundsel_4_5;
  wire roundsel_3_6;
  wire roundsel_2_6;
  wire roundsel_2_7;
  wire roundsel_2_8;
  wire roundsel_3_7;
  wire roundsel_3_8;
  wire roundsel_1_7;
  wire roundsel_1_8;
  wire roundsel_1_9;
  wire roundsel_3_5;
  wire roundsel_2_5;
  wire roundsel_2_10;
  wire roundsel_1_14;
  wire roundsel_4_6;
  wire roundsel_4_7;
  wire roundsel_4_8;
  wire roundsel_4_9;
  wire roundsel_3_10;
  wire roundsel_3_11;
  wire roundsel_3_12;
  wire roundsel_3_13;
  wire roundsel_3_14;
  wire roundsel_3_15;
  wire roundsel_1_15;
  wire roundsel_1_16;
  wire roundsel_1_17;
  wire roundsel_1_18;
  wire roundsel_1_19;
  wire roundsel_2_11;
  wire roundsel_2_12;
  wire roundsel_2_13;
  wire roundsel_1_20;
  wire roundsel_1_21;
  wire roundsel_1_22;
  wire roundsel_3_16;
  wire N5620;
  wire N5621;
  wire N5622;
  wire N5623;
  wire N5624;
  wire N5625;
  wire N5626;
  wire N5627;
  wire N5628;
  wire N5629;
  wire N5630;
  wire N5631;
  wire N5632;
  wire N5633;
  wire N5634;
  wire N5635;
  wire N5636;
  wire N5637;
  wire N5638;
  wire N5639;
  wire N5640;
  wire N5641;
  wire N5642;
  wire N5643;
  wire N5644;
  wire N5645;
  wire N5646;
  wire N5647;
  wire N5648;
  wire N5649;
  wire N5650;
  wire N5651;
  wire N5652;
  wire N5653;
  wire N5654;
  wire N5655;
  wire N5656;
  wire N5657;
  wire N5658;
  wire N5659;
  wire N5660;
  wire N5661;
  wire N5662;
  wire N5663;
  wire N5664;
  wire N5665;
  wire N5666;
  wire N5667;
  wire N5668;
  wire N5669;
  wire N5670;
  wire N5671;
  wire N5672;
  wire N5673;
  wire N5674;
  wire N5675;
  wire N5676;
  wire N5677;
  wire N5678;
  wire N5679;
  wire N5680;
  wire N5681;
  wire N5682;
  wire N5683;
  wire N5684;
  wire N5685;
  wire N5686;
  wire N5687;
  wire N5688;
  wire N5689;
  wire N5690;
  wire N5691;
  wire N5692;
  wire N5693;
  wire N5694;
  wire N5695;
  wire N5696;
  wire N5697;
  wire N5698;
  wire N5699;
  wire N5700;
  wire N5701;
  wire N5702;
  wire N5703;
  wire N5704;
  wire N5705;
  wire N5706;
  wire N5707;
  wire N5708;
  wire N5709;
  wire N5710;
  wire N5711;
  wire N5712;
  wire N5713;
  wire N5714;
  wire N5715;
  wire N5716;
  wire N5717;
  wire N5718;
  wire N5719;
  wire N5720;
  wire N5721;
  wire N5722;
  wire N5723;
  wire N5724;
  wire N5725;
  wire N5726;
  wire N5727;
  wire N5728;
  wire N5729;
  wire N5730;
  wire N5731;
  wire N5732;
  wire N5733;
  wire N5734;
  wire N5735;
  wire N5736;
  wire N5737;
  wire N5738;
  wire N5739;
  wire N5740;
  wire N5741;
  wire N5742;
  wire N5743;
  wire N5744;
  wire N5745;
  wire N5746;
  wire N5747;
  wire N5748;
  wire N5749;
  wire N5750;
  wire N5751;
  wire N5752;
  wire N5753;
  wire N5754;
  wire N5755;
  wire N5756;
  wire N5757;
  wire N5758;
  wire N5759;
  wire N5760;
  wire N5761;
  wire N5762;
  wire N5763;
  wire N5764;
  wire N5765;
  wire N5766;
  wire N5767;
  wire N5768;
  wire N5769;
  wire N5770;
  wire N5771;
  wire N5772;
  wire N5773;
  wire N5774;
  wire N5775;
  wire N5776;
  wire N5777;
  wire N5778;
  wire N5779;
  wire N5780;
  wire N5781;
  wire N5782;
  wire N5783;
  wire N5784;
  wire N5785;
  wire N5786;
  wire N5787;
  wire N5788;
  wire N5789;
  wire N5790;
  wire N5791;
  wire N5792;
  wire N5793;
  wire N5794;
  wire N5795;
  wire N5796;
  wire N5797;
  wire N5798;
  wire N5799;
  wire N5800;
  wire N5801;
  wire N5802;
  wire N5803;
  wire N5804;
  wire N5805;
  wire N5806;
  wire N5807;
  wire N5808;
  wire N5809;
  wire N5810;
  wire N5811;
  wire N5812;
  wire N5813;
  wire N5814;
  wire N5815;
  wire N5816;
  wire N5817;
  wire N5818;
  wire N5819;
  wire N5820;
  wire N5821;
  wire N5822;
  wire N5823;
  wire N5824;
  wire N5825;
  wire N5826;
  wire N5827;
  wire N5828;
  wire N5829;
  wire N5830;
  wire N5831;
  wire N5832;
  wire N5833;
  wire N5834;
  wire N5835;
  wire N5836;
  wire N5837;
  wire N5838;
  wire N5839;
  wire N5840;
  wire N5841;
  wire N5842;
  wire N5843;
  wire N5844;
  wire N5845;
  wire N5846;
  wire N5847;
  wire N5848;
  wire N5849;
  wire N5850;
  wire N5851;
  wire N5852;
  wire N5853;
  wire N5854;
  wire N5855;
  wire N5856;
  wire N5857;
  wire N5858;
  wire N5859;
  wire N5860;
  wire N5861;
  wire N5862;
  wire N5863;
  wire N5864;
  wire N5865;
  wire N5866;
  wire N5867;
  wire N5868;
  wire N5869;
  wire N5870;
  wire N5871;
  wire N5872;
  wire N5873;
  wire N5874;
  wire N5875;
  wire N5876;
  wire N5877;
  wire N5878;
  wire N5879;
  wire N5880;
  wire N5881;
  wire N5882;
  wire N5883;
  wire N5884;
  wire N5885;
  wire N5886;
  wire N5887;
  wire N5888;
  wire N5889;
  wire N5890;
  wire N5891;
  wire N5892;
  wire N5893;
  wire N5894;
  wire N5895;
  wire N5896;
  wire N5898;
  wire N5899;
  wire N5900;
  wire N5901;
  wire N5902;
  wire N5903;
  wire N5904;
  wire N5905;
  wire N5906;
  wire N5907;
  wire N5908;
  wire N5909;
  wire N5910;
  wire N5911;
  wire N5912;
  wire N5913;
  wire N5914;
  wire N5915;
  wire N5916;
  wire N5917;
  wire N5918;
  wire N5919;
  wire N5920;
  wire N5921;
  wire N5922;
  wire N5923;
  wire N5924;
  wire N5925;
  wire N5926;
  wire N5927;
  wire N5928;
  wire N5929;
  wire N5930;
  wire N5931;
  wire N5932;
  wire N5933;
  wire N5934;
  wire N5935;
  wire N5936;
  wire N5937;
  wire N5938;
  wire N5939;
  wire N5940;
  wire \key2<7>12_F/O ;
  wire \_n0013<6>22/O ;
  wire \key2<22>110_SW01_G/O ;
  wire \_n0013<8>22/O ;
  wire \_n0013<13>20/O ;
  wire \_n0013<10>22/O ;
  wire \key2<4>110_SW01_G/O ;
  wire \_n0013<0>22/O ;
  wire \_n0013<2>22/O ;
  wire \_n0013<7>20/O ;
  wire \_n0013<4>22/O ;
  wire \key2<3>1181_G/O ;
  wire \_n0013<63>22/O ;
  wire \_n0013<32>21/O ;
  wire \_n0013<61>22/O ;
  wire \key2<32>271_G/O ;
  wire \_n0013<59>22/O ;
  wire \_n0013<48>5/O ;
  wire \_n0013<57>22/O ;
  wire \_n0013<55>22/O ;
  wire \_n0013<53>22/O ;
  wire \_n0013<57>22_SW0/O ;
  wire \_n0013<51>22/O ;
  wire \_n0013<8>22_SW0/O ;
  wire \_n0013<49>22/O ;
  wire \key2<47>110_SW01_G/O ;
  wire \_n0013<47>22/O ;
  wire \_n0013<45>17/O ;
  wire \key2<28>1191_G/O ;
  wire \_n0013<43>22/O ;
  wire \_n0013<41>22/O ;
  wire \_n0013<39>22/O ;
  wire \_n0013<37>22/O ;
  wire \_n0013<35>22/O ;
  wire \_n0013<34>5/O ;
  wire \_n0013<33>22/O ;
  wire \_n0013<48>14/O ;
  wire \_n0013<30>22/O ;
  wire \_n0013<28>22/O ;
  wire \key2<25>961_G/O ;
  wire \_n0013<26>22/O ;
  wire \_n0013<24>22/O ;
  wire \key2<37>961_G/O ;
  wire \_n0013<22>22/O ;
  wire \_n0013<20>22/O ;
  wire \_n0013<17>20/O ;
  wire \_n0013<18>17/O ;
  wire \_n0013<13>20_SW1/O ;
  wire \_n0013<16>22/O ;
  wire \key2<38>961_G/O ;
  wire \_n0013<14>22/O ;
  wire \_n0013<12>22/O ;
  wire \key2<3>133_SW01_G/O ;
  wire \_n0013<14>22_SW0/O ;
  wire \key2<25>110_SW0/O ;
  wire \key2<25>12_SW0_G/O ;
  wire \key2<21>1191_G/O ;
  wire \key2<33>961_G/O ;
  wire \_n0013<1>20_SW0/O ;
  wire \key2<13>110_SW0/O ;
  wire \roundsel<2>_mmx_out271_G/O ;
  wire \key2<21>133_SW0/O ;
  wire \key2<27>156_SW0/O ;
  wire \key2<37>110_SW0/O ;
  wire \key2<28>133_SW0/O ;
  wire \key2<22>961_G/O ;
  wire \key2<45>133_SW0/O ;
  wire \_n0013<29>20_SW0_SW0/O ;
  wire \key2<43>110_SW0/O ;
  wire \key2<32>12_G/O ;
  wire \roundsel<1>_mmx_out621/O ;
  wire \roundsel<1>_mmx_out751/O ;
  wire \roundsel<2>_mmx_out71_G/O ;
  wire \key2<29>133_SW01_G/O ;
  wire \key2<41>961_G/O ;
  wire \key2<19>761_G/O ;
  wire \roundsel<2>_mmx_out111_G/O ;
  wire \key2<39>761_G/O ;
  wire \_n0013<11>20/O ;
  wire \_n0013<31>20_SW0_SW0/O ;
  wire \key2<31>761_G/O ;
  wire \key2<4>961_G/O ;
  wire \_n0013<23>20/O ;
  wire \key2<47>961_G/O ;
  wire \key2<17>25_SW0/O ;
  wire \key2<44>110_SW01_G/O ;
  wire \key2<34>110_SW01_G/O ;
  wire \key2<43>961_G/O ;
  wire \c1/Mxor_X_Result<7>11_G/O ;
  wire \key2<35>761_G/O ;
  wire \key2<45>471_G/O ;
  wire \_n0013<3>20_SW0/O ;
  wire \key2<6>110_SW01_G/O ;
  wire \key2<34>961_G/O ;
  wire \key2<6>961_G/O ;
  wire \key2<35>90_SW01_G/O ;
  wire \key2<30>1181_G/O ;
  wire \key2<17>471_G/O ;
  wire \key2<18>961_G/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_321/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_341/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_381/O ;
  wire \c1/u5/Mrom_dout_inst_mux_f5_18/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_401/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_421/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_441/O ;
  wire \c1/u5/Mrom_dout_inst_lut4_461/O ;
  wire \c1/Mxor_OUTR_Result<16>11_G/O ;
  wire \key2<42>110_SW01_G/O ;
  wire \key2<40>90_SW01_G/O ;
  wire \key2<21>471_G/O ;
  wire \key2<24>1181_G/O ;
  wire \key2<48>961_G/O ;
  wire \key2<36>1181_G/O ;
  wire \key2<23>1181_G/O ;
  wire \key2<48>110_SW01_G/O ;
  wire \c1/Mxor_X_Result<0>11_G/O ;
  wire \key2<1>271_G/O ;
  wire \key2<44>961_G/O ;
  wire \key2<18>110_SW01_G/O ;
  wire \key2<36>133_SW01_G/O ;
  wire \key2<16>271_G/O ;
  wire \c1/Mxor_X_Result<25>11_G/O ;
  wire \key2<14>1181_G/O ;
  wire \key2<12>761_G/O ;
  wire \c1/u3/Mrom_dout_inst_lut4_781/O ;
  wire \key2<8>61_G/O ;
  wire \c1/u3/Mrom_dout_inst_mux_f5_38/O ;
  wire \key2<13>961_G/O ;
  wire \key2<19>90_SW0/O ;
  wire \c1/Mxor_OUTR_Result<2>11_G/O ;
  wire \key2<9>471_G/O ;
  wire \c1/Mxor_OUTR_Result<1>11_G/O ;
  wire \c1/Mxor_OUTR_Result<9>11_G/O ;
  wire \key2<38>110_SW01_G/O ;
  wire \c1/Mxor_OUTR_Result<15>11_G/O ;
  wire \c1/Mxor_OUTR_Result<8>11_G/O ;
  wire \key2<41>110_SW01_G/O ;
  wire \c1/Mxor_OUTR_Result<26>11_G/O ;
  wire \c1/Mxor_OUTR_Result<29>11_G/O ;
  wire \c1/Mxor_OUTR_Result<22>11_G/O ;
  wire \c1/u1/Mrom_dout_inst_lut4_1141/O ;
  wire \c1/u1/Mrom_dout_inst_mux_f5_56/O ;
  wire \c1/u1/Mrom_dout_inst_lut4_1161/O ;
  wire \c1/u1/Mrom_dout_inst_lut4_1181/O ;
  wire \c1/u1/Mrom_dout_inst_lut4_1201/O ;
  wire \c1/u1/Mrom_dout_inst_lut4_1221/O ;
  wire \c1/u1/Mrom_dout_inst_mux_f5_62_SW1/O ;
  wire \c1/u1/Mrom_dout_inst_mux_f5_63_SW1/O ;
  wire \c1/Mxor_OUTR_Result<12>11_G/O ;
  wire \key2<12>90_SW0_G/O ;
  wire \c1/Mxor_OUTR_Result<6>11_G/O ;
  wire \key2<46>471_G/O ;
  wire \_n0013<48>21/O ;
  wire \_n0013<28>22_SW0/O ;
  wire \c1/Mxor_OUTR_Result<27>11_G/O ;
  wire \c1/Mxor_OUTR_Result<11>11_G/O ;
  wire \c1/Mxor_OUTR_Result<23>11_G/O ;
  wire \_n0013<42>5/O ;
  wire \_n0013<47>22_SW0/O ;
  wire \c1/Mxor_OUTR_Result<10>11_G/O ;
  wire \key2<8>271_G/O ;
  wire \_n0013<46>5/O ;
  wire \_n0013<34>14/O ;
  wire \_n0013<42>14/O ;
  wire \c1/Mxor_OUTR_Result<5>11_G/O ;
  wire \_n0013<42>21/O ;
  wire \_n0013<34>21/O ;
  wire \key2<40>761_G/O ;
  wire \_n0013<46>14/O ;
  wire \_n0013<30>1/O ;
  wire \_n0013<62>5/O ;
  wire \c1/Mxor_OUTR_Result<18>11_G/O ;
  wire \_n0013<46>21/O ;
  wire \c1/Mxor_OUTR_Result<0>11_G/O ;
  wire \_n0013<59>22_SW0/O ;
  wire \_n0013<2>22_SW0/O ;
  wire \_n0013<62>14/O ;
  wire \c1/Mxor_OUTR_Result<17>11_G/O ;
  wire \_n0013<62>21/O ;
  wire \_n0013<44>5/O ;
  wire \key2<2>961_G/O ;
  wire \_n0013<60>5/O ;
  wire \key2<26>271_G/O ;
  wire \_n0013<6>22_SW0/O ;
  wire \_n0013<44>14/O ;
  wire \key2<29>1181_G/O ;
  wire \key2<15>12/O ;
  wire \key2<15>1191_G/O ;
  wire \_n0013<60>14/O ;
  wire \_n0013<44>21/O ;
  wire \key2<20>961_G/O ;
  wire \_n0013<60>21/O ;
  wire \key2<37>271_G/O ;
  wire \key2<11>110_SW01_G/O ;
  wire \key2<25>271_G/O ;
  wire \key2<11>961_G/O ;
  wire \_n0013<58>5/O ;
  wire \_n0013<40>5/O ;
  wire \key2<39>90_SW01_G/O ;
  wire \_n0013<61>22_SW0/O ;
  wire \_n0013<51>22_SW0/O ;
  wire \_n0013<58>14/O ;
  wire \_n0013<58>21/O ;
  wire \_n0013<40>14/O ;
  wire \_n0013<0>22_SW0/O ;
  wire \_n0013<40>21/O ;
  wire \key2<23>133_SW01_G/O ;
  wire \key2<30>133_SW01_G/O ;
  wire \key2<46>1191_G/O ;
  wire \_n0013<54>5/O ;
  wire \_n0013<37>22_SW0/O ;
  wire \key2<13>271_G/O ;
  wire \key2<42>961_G/O ;
  wire \_n0013<38>5/O ;
  wire \_n0013<54>14/O ;
  wire \_n0013<9>20_SW0_SW0_SW0_SW0/O ;
  wire \key2<10>961_G/O ;
  wire \_n0013<54>21/O ;
  wire \key2<15>471_G/O ;
  wire \key2<9>1191_G/O ;
  wire \key2<27>471_G/O ;
  wire \_n0013<38>14/O ;
  wire \_n0013<56>5/O ;
  wire \c1/Mxor_X_Result<31>11_G/O ;
  wire \_n0013<39>12/O ;
  wire \_n0013<38>21/O ;
  wire \key2<24>133_SW01_G/O ;
  wire \_n0013<56>14/O ;
  wire \key2<27>1411_G/O ;
  wire \key2<10>110_SW01_G/O ;
  wire \_n0013<56>21/O ;
  wire \key2<2>110_SW01_G/O ;
  wire \key2<5>110_SW01_G/O ;
  wire \_n0013<36>5/O ;
  wire \_n0013<10>22_SW0/O ;
  wire \_n0013<18>17_SW0/O ;
  wire \_n0013<52>5/O ;
  wire \key2<7>761_G/O ;
  wire \key2<33>110_SW01_G/O ;
  wire \key2<45>1191_G/O ;
  wire \key2<5>961_G/O ;
  wire \key2<14>133_SW01_G/O ;
  wire \_n0013<36>14/O ;
  wire \_n0013<41>22_SW0/O ;
  wire \_n0013<52>14/O ;
  wire \key2<43>271_G/O ;
  wire \_n0013<55>22_SW0/O ;
  wire \_n0013<36>21/O ;
  wire \_n0013<52>21/O ;
  wire \c1/Mxor_X_Result<15>11_G/O ;
  wire \key2<28>471_G/O ;
  wire \key2<17>1191_G/O ;
  wire \key2<20>110_SW01_G/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_291_G/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_281_G/O ;
  wire \_n0013<50>5/O ;
  wire \_n0013<32>5/O ;
  wire \roundsel<2>_mmx_out331_G/O ;
  wire \_n0013<50>14/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_251_G/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_241_G/O ;
  wire \_n0013<50>21/O ;
  wire \c1/u6/Mrom_dout_inst_mux_f5_111_G/O ;
  wire \_n0013<32>14/O ;
  wire \Ker020_SW0/O ;
  wire \_n0013<26>22_SW0/O ;
  wire \_n0013<7>20_SW0/O ;
  wire \c1/u6/Mrom_dout_inst_mux_f5_101_G/O ;
  wire \_n0013<15>20/O ;
  wire \c1/Mxor_OUTR_Result<25>11_G/O ;
  wire \_n0013<27>20_SW0/O ;
  wire \roundsel<2>_mmx_out241_G/O ;
  wire \key2<31>15_G/O ;
  wire \key2<9>12/O ;
  wire \_n0013<3>20/O ;
  wire \key2<46>12/O ;
  wire \key2<26>12_G/O ;
  wire \_n0013<11>20_SW0/O ;
  wire \_n0013<1>20/O ;
  wire \_n0013<19>20/O ;
  wire \_n0013<9>20/O ;
  wire \_n0013<19>20_SW0/O ;
  wire \key2<8>12_G/O ;
  wire \_n0013<21>20/O ;
  wire \_n0013<21>20_SW0/O ;
  wire \_n0013<23>20_SW0/O ;
  wire \_n0013<25>20/O ;
  wire \key2<37>12_SW0_G/O ;
  wire \_n0013<15>20_SW0/O ;
  wire \_n0013<29>20/O ;
  wire \_n0013<20>22_SW0/O ;
  wire \_n0013<16>22_SW0/O ;
  wire \_n0013<17>20_SW0/O ;
  wire \_n0013<5>20_SW0/O ;
  wire \_n0013<27>20/O ;
  wire \key2<43>12_SW0_G/O ;
  wire \_n0013<25>20_SW0/O ;
  wire \_n0013<5>20/O ;
  wire \_n0013<12>22_SW0/O ;
  wire \key2<13>12_SW0_G/O ;
  wire \_n0013<22>22_SW0/O ;
  wire \_n0013<31>20/O ;
  wire \Ker039_1/O ;
  wire \key2<7>15_G/O ;
  wire \key2<26>61_G/O ;
  wire \key2<31>12_G/O ;
  wire \key2<7>12_G/O ;
  wire \key2<22>110_SW01_F/O ;
  wire \key2<4>110_SW01_F/O ;
  wire \key2<3>1181_F/O ;
  wire \key2<32>271_F/O ;
  wire \key2<47>110_SW01_F/O ;
  wire \key2<28>1191_F/O ;
  wire \key2<25>961_F/O ;
  wire \key2<37>961_F/O ;
  wire \key2<38>961_F/O ;
  wire \key2<3>133_SW01_F/O ;
  wire \key2<25>12_SW0_F/O ;
  wire \key2<21>1191_F/O ;
  wire \key2<33>961_F/O ;
  wire \roundsel<2>_mmx_out271_F/O ;
  wire \key2<22>961_F/O ;
  wire \key2<32>12_F/O ;
  wire \roundsel<2>_mmx_out71_F/O ;
  wire \key2<29>133_SW01_F/O ;
  wire \key2<41>961_F/O ;
  wire \key2<19>761_F/O ;
  wire \roundsel<2>_mmx_out111_F/O ;
  wire \key2<39>761_F/O ;
  wire \key2<31>761_F/O ;
  wire \key2<4>961_F/O ;
  wire \key2<47>961_F/O ;
  wire \key2<44>110_SW01_F/O ;
  wire \key2<34>110_SW01_F/O ;
  wire \key2<43>961_F/O ;
  wire \c1/Mxor_X_Result<7>11_F/O ;
  wire \key2<35>761_F/O ;
  wire \key2<45>471_F/O ;
  wire \key2<6>110_SW01_F/O ;
  wire \key2<34>961_F/O ;
  wire \key2<6>961_F/O ;
  wire \key2<35>90_SW01_F/O ;
  wire \key2<30>1181_F/O ;
  wire \key2<17>471_F/O ;
  wire \key2<18>961_F/O ;
  wire \c1/Mxor_OUTR_Result<16>11_F/O ;
  wire \key2<42>110_SW01_F/O ;
  wire \key2<40>90_SW01_F/O ;
  wire \key2<21>471_F/O ;
  wire \key2<24>1181_F/O ;
  wire \key2<48>961_F/O ;
  wire \key2<36>1181_F/O ;
  wire \key2<23>1181_F/O ;
  wire \key2<48>110_SW01_F/O ;
  wire \c1/Mxor_X_Result<0>11_F/O ;
  wire \key2<1>271_F/O ;
  wire \key2<44>961_F/O ;
  wire \key2<18>110_SW01_F/O ;
  wire \key2<36>133_SW01_F/O ;
  wire \key2<16>271_F/O ;
  wire \c1/Mxor_X_Result<25>11_F/O ;
  wire \key2<14>1181_F/O ;
  wire \key2<12>761_F/O ;
  wire \key2<8>61_F/O ;
  wire \key2<13>961_F/O ;
  wire \c1/Mxor_OUTR_Result<2>11_F/O ;
  wire \key2<9>471_F/O ;
  wire \c1/Mxor_OUTR_Result<1>11_F/O ;
  wire \c1/Mxor_OUTR_Result<9>11_F/O ;
  wire \key2<38>110_SW01_F/O ;
  wire \c1/Mxor_OUTR_Result<15>11_F/O ;
  wire \c1/Mxor_OUTR_Result<8>11_F/O ;
  wire \key2<41>110_SW01_F/O ;
  wire \c1/Mxor_OUTR_Result<26>11_F/O ;
  wire \c1/Mxor_OUTR_Result<29>11_F/O ;
  wire \c1/Mxor_OUTR_Result<22>11_F/O ;
  wire \c1/Mxor_OUTR_Result<12>11_F/O ;
  wire \key2<12>90_SW0_F/O ;
  wire \c1/Mxor_OUTR_Result<6>11_F/O ;
  wire \key2<46>471_F/O ;
  wire \c1/Mxor_OUTR_Result<27>11_F/O ;
  wire \c1/Mxor_OUTR_Result<11>11_F/O ;
  wire \c1/Mxor_OUTR_Result<23>11_F/O ;
  wire \c1/Mxor_OUTR_Result<10>11_F/O ;
  wire \key2<8>271_F/O ;
  wire \c1/Mxor_OUTR_Result<5>11_F/O ;
  wire \key2<40>761_F/O ;
  wire \c1/Mxor_OUTR_Result<18>11_F/O ;
  wire \c1/Mxor_OUTR_Result<0>11_F/O ;
  wire \c1/Mxor_OUTR_Result<17>11_F/O ;
  wire \key2<2>961_F/O ;
  wire \key2<26>271_F/O ;
  wire \key2<29>1181_F/O ;
  wire \key2<15>1191_F/O ;
  wire \key2<20>961_F/O ;
  wire \key2<37>271_F/O ;
  wire \key2<11>110_SW01_F/O ;
  wire \key2<25>271_F/O ;
  wire \key2<11>961_F/O ;
  wire \key2<39>90_SW01_F/O ;
  wire \key2<23>133_SW01_F/O ;
  wire \key2<30>133_SW01_F/O ;
  wire \key2<46>1191_F/O ;
  wire \key2<13>271_F/O ;
  wire \key2<42>961_F/O ;
  wire \key2<10>961_F/O ;
  wire \key2<15>471_F/O ;
  wire \key2<9>1191_F/O ;
  wire \key2<27>471_F/O ;
  wire \c1/Mxor_X_Result<31>11_F/O ;
  wire \key2<24>133_SW01_F/O ;
  wire \key2<27>1411_F/O ;
  wire \key2<10>110_SW01_F/O ;
  wire \key2<2>110_SW01_F/O ;
  wire \key2<5>110_SW01_F/O ;
  wire \key2<7>761_F/O ;
  wire \key2<33>110_SW01_F/O ;
  wire \key2<45>1191_F/O ;
  wire \key2<5>961_F/O ;
  wire \key2<14>133_SW01_F/O ;
  wire \key2<43>271_F/O ;
  wire \c1/Mxor_X_Result<15>11_F/O ;
  wire \key2<28>471_F/O ;
  wire \key2<17>1191_F/O ;
  wire \key2<20>110_SW01_F/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_291_F/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_281_F/O ;
  wire \roundsel<2>_mmx_out331_F/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_251_F/O ;
  wire \c1/u4/Mrom_dout_inst_mux_f5_241_F/O ;
  wire \c1/u6/Mrom_dout_inst_mux_f5_111_F/O ;
  wire \c1/u6/Mrom_dout_inst_mux_f5_101_F/O ;
  wire \c1/Mxor_OUTR_Result<25>11_F/O ;
  wire \roundsel<2>_mmx_out241_F/O ;
  wire \key2<31>15_F/O ;
  wire \key2<26>12_F/O ;
  wire \key2<8>12_F/O ;
  wire \key2<37>12_SW0_F/O ;
  wire \key2<43>12_SW0_F/O ;
  wire \key2<13>12_SW0_F/O ;
  wire \key2<7>15_F/O ;
  wire \key2<26>61_F/O ;
  wire \key2<31>12_F/O ;
  wire \clk_BUFGP/IBUFG ;
  wire GSR = glbl.GSR;
  wire \dataout_1_OBUF.GTS.TRI ;
  wire GTS = glbl.GTS;
  wire \dataout_23_OBUF.GTS.TRI ;
  wire \dataout_4_OBUF.GTS.TRI ;
  wire \dataout_48_OBUF.GTS.TRI ;
  wire \dataout_43_OBUF.GTS.TRI ;
  wire \dataout_25_OBUF.GTS.TRI ;
  wire \dataout_49_OBUF.GTS.TRI ;
  wire \dataout_31_OBUF.GTS.TRI ;
  wire \dataout_24_OBUF.GTS.TRI ;
  wire \dataout_35_OBUF.GTS.TRI ;
  wire \dataout_33_OBUF.GTS.TRI ;
  wire \dataout_46_OBUF.GTS.TRI ;
  wire \dataout_26_OBUF.GTS.TRI ;
  wire \dataout_17_OBUF.GTS.TRI ;
  wire \dataout_45_OBUF.GTS.TRI ;
  wire \dataout_40_OBUF.GTS.TRI ;
  wire \dataout_42_OBUF.GTS.TRI ;
  wire \dataout_6_OBUF.GTS.TRI ;
  wire \dataout_3_OBUF.GTS.TRI ;
  wire \dataout_51_OBUF.GTS.TRI ;
  wire \dataout_28_OBUF.GTS.TRI ;
  wire \dataout_5_OBUF.GTS.TRI ;
  wire \dataout_37_OBUF.GTS.TRI ;
  wire \dataout_36_OBUF.GTS.TRI ;
  wire \dataout_30_OBUF.GTS.TRI ;
  wire \dataout_39_OBUF.GTS.TRI ;
  wire \dataout_32_OBUF.GTS.TRI ;
  wire \dataout_29_OBUF.GTS.TRI ;
  wire \dataout_27_OBUF.GTS.TRI ;
  wire \dataout_34_OBUF.GTS.TRI ;
  wire \dataout_47_OBUF.GTS.TRI ;
  wire \dataout_38_OBUF.GTS.TRI ;
  wire \dataout_41_OBUF.GTS.TRI ;
  wire \dataout_50_OBUF.GTS.TRI ;
  wire \dataout_44_OBUF.GTS.TRI ;
  wire \dataout_2_OBUF.GTS.TRI ;
  wire \ready_OBUF.GTS.TRI ;
  wire \dataout_15_OBUF.GTS.TRI ;
  wire \dataout_11_OBUF.GTS.TRI ;
  wire \dataout_14_OBUF.GTS.TRI ;
  wire \dataout_61_OBUF.GTS.TRI ;
  wire \dataout_7_OBUF.GTS.TRI ;
  wire \dataout_63_OBUF.GTS.TRI ;
  wire \dataout_64_OBUF.GTS.TRI ;
  wire \dataout_8_OBUF.GTS.TRI ;
  wire \dataout_52_OBUF.GTS.TRI ;
  wire \dataout_9_OBUF.GTS.TRI ;
  wire \dataout_56_OBUF.GTS.TRI ;
  wire \dataout_21_OBUF.GTS.TRI ;
  wire \dataout_62_OBUF.GTS.TRI ;
  wire \dataout_57_OBUF.GTS.TRI ;
  wire \dataout_19_OBUF.GTS.TRI ;
  wire \dataout_60_OBUF.GTS.TRI ;
  wire \dataout_58_OBUF.GTS.TRI ;
  wire \dataout_10_OBUF.GTS.TRI ;
  wire \dataout_55_OBUF.GTS.TRI ;
  wire \dataout_54_OBUF.GTS.TRI ;
  wire \dataout_12_OBUF.GTS.TRI ;
  wire \dataout_22_OBUF.GTS.TRI ;
  wire \dataout_16_OBUF.GTS.TRI ;
  wire \dataout_59_OBUF.GTS.TRI ;
  wire \dataout_13_OBUF.GTS.TRI ;
  wire \dataout_18_OBUF.GTS.TRI ;
  wire \dataout_53_OBUF.GTS.TRI ;
  wire \dataout_20_OBUF.GTS.TRI ;
  wire VCC;
  wire GND;
  wire \NlwInverterSignal_dataout_1_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_23_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_4_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_48_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_43_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_25_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_49_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_31_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_24_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_35_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_33_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_46_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_26_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_17_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_45_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_40_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_42_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_6_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_3_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_51_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_28_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_5_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_37_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_36_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_30_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_39_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_32_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_29_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_27_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_34_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_47_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_38_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_41_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_50_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_44_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_2_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_ready_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_15_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_11_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_14_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_61_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_7_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_63_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_64_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_8_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_52_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_9_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_56_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_21_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_62_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_57_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_19_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_60_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_58_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_10_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_55_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_54_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_12_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_22_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_16_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_59_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_13_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_18_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_53_OBUF.GTS.TRI/CTL ;
  wire \NlwInverterSignal_dataout_20_OBUF.GTS.TRI/CTL ;
  wire [0 : 0] _n0012;
  wire [64 : 1] data1;
  wire [63 : 0] _n0013;
  wire [4 : 1] roundsel;
  wire [32 : 1] cipherout2;
  wire [0 : 0] \Maddsub__n0017_Mxor_Result<3>_Xo ;
  wire [2 : 2] _n0032;
  defparam ready_0.INIT = 1'b0;
  X_SFF ready_0 (
    .I(N5011),
    .SRST(_n0032[2]),
    .SSET(state_FFd1),
    .CLK(clk_BUFGP),
    .O(ready_OBUF),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  X_ZERO XST_GND (
    .O(N1)
  );
  X_BUF key_42_IBUF_1 (
    .I(key[42]),
    .O(key_42_IBUF)
  );
  defparam _n00291.INIT = 4'h8;
  X_LUT2 _n00291 (
    .ADR0(state_FFd8),
    .ADR1(rst_IBUF),
    .O(_n0029)
  );
  defparam _n00301.INIT = 4'h8;
  X_LUT2 _n00301 (
    .ADR0(state_FFd3),
    .ADR1(rst_IBUF),
    .O(_n0030)
  );
  defparam \roundsel<1>_mmx_out861 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out861  (
    .ADR0(\key1[54] ),
    .ADR1(\key1[5] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out86 )
  );
  defparam _n00251.INIT = 4'hE;
  X_LUT2 _n00251 (
    .ADR0(state_FFd6),
    .ADR1(state_FFd5),
    .O(_n0025)
  );
  defparam data1_62.INIT = 1'b0;
  X_FF data1_62 (
    .I(_n0013[61]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[62]),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3.INIT = 1'b1;
  X_SFF roundsel_3 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel[3]),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam data1_60.INIT = 1'b0;
  X_FF data1_60 (
    .I(_n0013[59]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[60]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_61.INIT = 1'b0;
  X_FF data1_61 (
    .I(_n0013[60]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[61]),
    .SET(GND),
    .RST(GSR)
  );
  X_BUF datain_19_IBUF_2 (
    .I(datain[19]),
    .O(datain_19_IBUF)
  );
  defparam \roundsel<1>_mmx_out941 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out941  (
    .ADR0(\key1[14] ),
    .ADR1(\key1[63] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out94 )
  );
  X_BUF datain_21_IBUF_3 (
    .I(datain[21]),
    .O(datain_21_IBUF)
  );
  X_BUF datain_23_IBUF_4 (
    .I(datain[23]),
    .O(datain_23_IBUF)
  );
  X_BUF dataout_55_OBUF (
    .I(dataout_55),
    .O(\dataout_55_OBUF.GTS.TRI )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_63_SW0 .INIT = 16'h9621;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_63_SW0  (
    .ADR0(data1[29]),
    .ADR1(\c1/X[8] ),
    .ADR2(N5898),
    .ADR3(\c1/X[10] ),
    .O(N5183)
  );
  defparam state_FFd6_5.INIT = 1'b0;
  X_SFF state_FFd6_5 (
    .I(\state_FFd6-In ),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd6),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam state_FFd5_6.INIT = 1'b0;
  X_SFF state_FFd5_6 (
    .I(\state_FFd5-In ),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd5),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam _n00111.INIT = 8'hEA;
  X_LUT3 _n00111 (
    .ADR0(N234),
    .ADR1(_n0000),
    .ADR2(state_FFd4),
    .O(N5011)
  );
  defparam \_n0012<3>551 .INIT = 4'h8;
  X_LUT2 \_n0012<3>551  (
    .ADR0(rst_IBUF),
    .ADR1(CHOICE13),
    .O(N5008)
  );
  defparam data1_64.INIT = 1'b0;
  X_FF data1_64 (
    .I(_n0013[63]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[64]),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_64.INIT = 1'b0;
  X_FF key1_64 (
    .I(key_64_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[64] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_64_7.INIT = 1'b0;
  X_FF dataout_64_7 (
    .I(data1[64]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_64),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3_4.INIT = 1'b1;
  X_SFF roundsel_3_4 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_2),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  X_BUF datain_25_IBUF_8 (
    .I(datain[25]),
    .O(datain_25_IBUF)
  );
  X_BUF datain_58_IBUF_9 (
    .I(datain[58]),
    .O(datain_58_IBUF)
  );
  defparam \roundsel<1>_mmx_out841 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out841  (
    .ADR0(\key1[6] ),
    .ADR1(\key1[55] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out84 )
  );
  defparam roundsel_2.INIT = 1'b1;
  X_SFF roundsel_2 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel[2]),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  X_BUF dataout_58_OBUF (
    .I(dataout_58),
    .O(\dataout_58_OBUF.GTS.TRI )
  );
  defparam \key2<27>25_SW0 .INIT = 16'hF3F5;
  X_LUT4 \key2<27>25_SW0  (
    .ADR0(\key1[23] ),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_3_8),
    .ADR3(roundsel_12),
    .O(N5133)
  );
  defparam \_n0012<2>100_SW2 .INIT = 16'h77EF;
  X_LUT4 \_n0012<2>100_SW2  (
    .ADR0(roundsel[1]),
    .ADR1(roundsel[2]),
    .ADR2(state_FFd5),
    .ADR3(state_FFd6),
    .O(N5499)
  );
  defparam \_n0012<0>_G .INIT = 16'hF272;
  X_LUT4 \_n0012<0>_G  (
    .ADR0(rst_IBUF),
    .ADR1(roundsel[1]),
    .ADR2(flag_IBUF),
    .ADR3(state_FFd7),
    .O(N5633)
  );
  X_BUF key_5_IBUF_10 (
    .I(key[5]),
    .O(key_5_IBUF)
  );
  defparam \_n0013<28>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<28>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[33]),
    .ADR2(state_FFd8),
    .ADR3(datain_29_IBUF),
    .O(CHOICE831)
  );
  defparam \_n0013<57>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<57>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[10]),
    .ADR2(state_FFd8),
    .ADR3(datain_58_IBUF),
    .O(CHOICE713)
  );
  X_BUF ready_OBUF_11 (
    .I(ready_OBUF),
    .O(\ready_OBUF.GTS.TRI )
  );
  X_BUF dataout_21_OBUF (
    .I(dataout_21),
    .O(\dataout_21_OBUF.GTS.TRI )
  );
  X_BUF dataout_60_OBUF (
    .I(dataout_60),
    .O(\dataout_60_OBUF.GTS.TRI )
  );
  X_BUF key_48_IBUF_12 (
    .I(key[48]),
    .O(key_48_IBUF)
  );
  defparam \_n0013<13>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<13>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[45]),
    .ADR2(state_FFd8),
    .ADR3(datain_14_IBUF),
    .O(CHOICE2017)
  );
  defparam data1_63.INIT = 1'b0;
  X_FF data1_63 (
    .I(_n0013[62]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[63]),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1.INIT = 1'b0;
  X_FF roundsel_1 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel[1]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \_n0012<2>1271 .INIT = 4'h8;
  X_LUT2 \_n0012<2>1271  (
    .ADR0(rst_IBUF),
    .ADR1(CHOICE230),
    .O(N5010)
  );
  defparam dataout_1_13.INIT = 1'b0;
  X_FF dataout_1_13 (
    .I(data1[1]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_1),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_2_14.INIT = 1'b0;
  X_FF dataout_2_14 (
    .I(data1[2]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_2),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_3_15.INIT = 1'b0;
  X_FF dataout_3_15 (
    .I(data1[3]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_3),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_4_16.INIT = 1'b0;
  X_FF dataout_4_16 (
    .I(data1[4]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_4),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_5_17.INIT = 1'b0;
  X_FF dataout_5_17 (
    .I(data1[5]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_5),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_6_18.INIT = 1'b0;
  X_FF dataout_6_18 (
    .I(data1[6]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_6),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_7_19.INIT = 1'b0;
  X_FF dataout_7_19 (
    .I(data1[7]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_7),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_8_20.INIT = 1'b0;
  X_FF dataout_8_20 (
    .I(data1[8]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_8),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_9_21.INIT = 1'b0;
  X_FF dataout_9_21 (
    .I(data1[9]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_9),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_10_22.INIT = 1'b0;
  X_FF dataout_10_22 (
    .I(data1[10]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_10),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_11_23.INIT = 1'b0;
  X_FF dataout_11_23 (
    .I(data1[11]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_11),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_12_24.INIT = 1'b0;
  X_FF dataout_12_24 (
    .I(data1[12]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_12),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_13_25.INIT = 1'b0;
  X_FF dataout_13_25 (
    .I(data1[13]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_13),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_14_26.INIT = 1'b0;
  X_FF dataout_14_26 (
    .I(data1[14]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_14),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_15_27.INIT = 1'b0;
  X_FF dataout_15_27 (
    .I(data1[15]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_15),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_16_28.INIT = 1'b0;
  X_FF dataout_16_28 (
    .I(data1[16]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_16),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_17_29.INIT = 1'b0;
  X_FF dataout_17_29 (
    .I(data1[17]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_17),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_18_30.INIT = 1'b0;
  X_FF dataout_18_30 (
    .I(data1[18]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_18),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_19_31.INIT = 1'b0;
  X_FF dataout_19_31 (
    .I(data1[19]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_19),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_20_32.INIT = 1'b0;
  X_FF dataout_20_32 (
    .I(data1[20]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_20),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_21_33.INIT = 1'b0;
  X_FF dataout_21_33 (
    .I(data1[21]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_21),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_22_34.INIT = 1'b0;
  X_FF dataout_22_34 (
    .I(data1[22]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_22),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_23_35.INIT = 1'b0;
  X_FF dataout_23_35 (
    .I(data1[23]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_23),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_24_36.INIT = 1'b0;
  X_FF dataout_24_36 (
    .I(data1[24]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_24),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_25_37.INIT = 1'b0;
  X_FF dataout_25_37 (
    .I(data1[25]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_25),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_26_38.INIT = 1'b0;
  X_FF dataout_26_38 (
    .I(data1[26]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_26),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_27_39.INIT = 1'b0;
  X_FF dataout_27_39 (
    .I(data1[27]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_27),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_28_40.INIT = 1'b0;
  X_FF dataout_28_40 (
    .I(data1[28]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_28),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_29_41.INIT = 1'b0;
  X_FF dataout_29_41 (
    .I(data1[29]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_29),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_30_42.INIT = 1'b0;
  X_FF dataout_30_42 (
    .I(data1[30]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_30),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_31_43.INIT = 1'b0;
  X_FF dataout_31_43 (
    .I(data1[31]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_31),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_32_44.INIT = 1'b0;
  X_FF dataout_32_44 (
    .I(data1[32]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_32),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_33_45.INIT = 1'b0;
  X_FF dataout_33_45 (
    .I(data1[33]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_33),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_34_46.INIT = 1'b0;
  X_FF dataout_34_46 (
    .I(data1[34]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_34),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_35_47.INIT = 1'b0;
  X_FF dataout_35_47 (
    .I(data1[35]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_35),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_36_48.INIT = 1'b0;
  X_FF dataout_36_48 (
    .I(data1[36]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_36),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_37_49.INIT = 1'b0;
  X_FF dataout_37_49 (
    .I(data1[37]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_37),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_38_50.INIT = 1'b0;
  X_FF dataout_38_50 (
    .I(data1[38]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_38),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_39_51.INIT = 1'b0;
  X_FF dataout_39_51 (
    .I(data1[39]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_39),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_40_52.INIT = 1'b0;
  X_FF dataout_40_52 (
    .I(data1[40]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_40),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_41_53.INIT = 1'b0;
  X_FF dataout_41_53 (
    .I(data1[41]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_41),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_42_54.INIT = 1'b0;
  X_FF dataout_42_54 (
    .I(data1[42]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_42),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_43_55.INIT = 1'b0;
  X_FF dataout_43_55 (
    .I(data1[43]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_43),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_44_56.INIT = 1'b0;
  X_FF dataout_44_56 (
    .I(data1[44]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_44),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_45_57.INIT = 1'b0;
  X_FF dataout_45_57 (
    .I(data1[45]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_45),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_46_58.INIT = 1'b0;
  X_FF dataout_46_58 (
    .I(data1[46]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_46),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_47_59.INIT = 1'b0;
  X_FF dataout_47_59 (
    .I(data1[47]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_47),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_48_60.INIT = 1'b0;
  X_FF dataout_48_60 (
    .I(data1[48]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_48),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_49_61.INIT = 1'b0;
  X_FF dataout_49_61 (
    .I(data1[49]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_49),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_50_62.INIT = 1'b0;
  X_FF dataout_50_62 (
    .I(data1[50]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_50),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_51_63.INIT = 1'b0;
  X_FF dataout_51_63 (
    .I(data1[51]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_51),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_52_64.INIT = 1'b0;
  X_FF dataout_52_64 (
    .I(data1[52]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_52),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_53_65.INIT = 1'b0;
  X_FF dataout_53_65 (
    .I(data1[53]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_53),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_54_66.INIT = 1'b0;
  X_FF dataout_54_66 (
    .I(data1[54]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_54),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_55_67.INIT = 1'b0;
  X_FF dataout_55_67 (
    .I(data1[55]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_55),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_56_68.INIT = 1'b0;
  X_FF dataout_56_68 (
    .I(data1[56]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_56),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_57_69.INIT = 1'b0;
  X_FF dataout_57_69 (
    .I(data1[57]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_57),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_58_70.INIT = 1'b0;
  X_FF dataout_58_70 (
    .I(data1[58]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_58),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_59_71.INIT = 1'b0;
  X_FF dataout_59_71 (
    .I(data1[59]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_59),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_60_72.INIT = 1'b0;
  X_FF dataout_60_72 (
    .I(data1[60]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_60),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_61_73.INIT = 1'b0;
  X_FF dataout_61_73 (
    .I(data1[61]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_61),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_62_74.INIT = 1'b0;
  X_FF dataout_62_74 (
    .I(data1[62]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_62),
    .SET(GND),
    .RST(GSR)
  );
  defparam dataout_63_75.INIT = 1'b0;
  X_FF dataout_63_75 (
    .I(data1[63]),
    .CE(_n0030),
    .CLK(clk_BUFGP),
    .O(dataout_63),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd2_76.INIT = 1'b0;
  X_SFF state_FFd2_76 (
    .I(state_FFd5),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd2),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam key1_2.INIT = 1'b0;
  X_FF key1_2 (
    .I(key_2_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[2] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_3.INIT = 1'b0;
  X_FF key1_3 (
    .I(key_3_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[3] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_4.INIT = 1'b0;
  X_FF key1_4 (
    .I(key_4_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[4] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_5.INIT = 1'b0;
  X_FF key1_5 (
    .I(key_5_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[5] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_6.INIT = 1'b0;
  X_FF key1_6 (
    .I(key_6_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[6] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_7.INIT = 1'b0;
  X_FF key1_7 (
    .I(key_7_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[7] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_8.INIT = 1'b0;
  X_FF key1_8 (
    .I(key_8_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[8] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd1_77.INIT = 1'b0;
  X_SFF state_FFd1_77 (
    .I(state_FFd3),
    .SRST(_n0032[2]),
    .SSET(state_FFd1),
    .CLK(clk_BUFGP),
    .O(state_FFd1),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_10.INIT = 1'b0;
  X_FF key1_10 (
    .I(key_10_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[10] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_11.INIT = 1'b0;
  X_FF key1_11 (
    .I(key_11_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[11] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_12.INIT = 1'b0;
  X_FF key1_12 (
    .I(key_12_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[12] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_13.INIT = 1'b0;
  X_FF key1_13 (
    .I(key_13_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[13] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_14.INIT = 1'b0;
  X_FF key1_14 (
    .I(key_14_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[14] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_15.INIT = 1'b0;
  X_FF key1_15 (
    .I(key_15_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[15] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_16.INIT = 1'b0;
  X_FF key1_16 (
    .I(key_16_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[16] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd3_78.INIT = 1'b0;
  X_SFF state_FFd3_78 (
    .I(N5899),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd3),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam key1_18.INIT = 1'b0;
  X_FF key1_18 (
    .I(key_18_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[18] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_19.INIT = 1'b0;
  X_FF key1_19 (
    .I(key_19_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[19] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_20.INIT = 1'b0;
  X_FF key1_20 (
    .I(key_20_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[20] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_21.INIT = 1'b0;
  X_FF key1_21 (
    .I(key_21_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[21] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_22.INIT = 1'b0;
  X_FF key1_22 (
    .I(key_22_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[22] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_23.INIT = 1'b0;
  X_FF key1_23 (
    .I(key_23_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[23] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_24.INIT = 1'b0;
  X_FF key1_24 (
    .I(key_24_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[24] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd8_79.INIT = 1'b1;
  X_SFF state_FFd8_79 (
    .I(N1),
    .SSET(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd8),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam key1_26.INIT = 1'b0;
  X_FF key1_26 (
    .I(key_26_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[26] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_27.INIT = 1'b0;
  X_FF key1_27 (
    .I(key_27_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[27] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_28.INIT = 1'b0;
  X_FF key1_28 (
    .I(key_28_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[28] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_29.INIT = 1'b0;
  X_FF key1_29 (
    .I(key_29_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[29] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_30.INIT = 1'b0;
  X_FF key1_30 (
    .I(key_30_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[30] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_31.INIT = 1'b0;
  X_FF key1_31 (
    .I(key_31_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[31] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_32.INIT = 1'b0;
  X_FF key1_32 (
    .I(key_32_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[32] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \state_FFd6-In1 .INIT = 16'h4F44;
  X_LUT4 \state_FFd6-In1  (
    .ADR0(flag_IBUF),
    .ADR1(state_FFd7),
    .ADR2(_n0000),
    .ADR3(state_FFd4),
    .O(\state_FFd6-In )
  );
  defparam key1_34.INIT = 1'b0;
  X_FF key1_34 (
    .I(key_34_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[34] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_35.INIT = 1'b0;
  X_FF key1_35 (
    .I(key_35_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[35] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_36.INIT = 1'b0;
  X_FF key1_36 (
    .I(key_36_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[36] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_37.INIT = 1'b0;
  X_FF key1_37 (
    .I(key_37_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[37] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_38.INIT = 1'b0;
  X_FF key1_38 (
    .I(key_38_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[38] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_39.INIT = 1'b0;
  X_FF key1_39 (
    .I(key_39_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[39] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_40.INIT = 1'b0;
  X_FF key1_40 (
    .I(key_40_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[40] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \state_FFd5-In1 .INIT = 16'hF444;
  X_LUT4 \state_FFd5-In1  (
    .ADR0(_n0001),
    .ADR1(state_FFd2),
    .ADR2(flag_IBUF),
    .ADR3(state_FFd7),
    .O(\state_FFd5-In )
  );
  defparam key1_42.INIT = 1'b0;
  X_FF key1_42 (
    .I(key_42_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[42] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_43.INIT = 1'b0;
  X_FF key1_43 (
    .I(key_43_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[43] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_44.INIT = 1'b0;
  X_FF key1_44 (
    .I(key_44_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[44] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_45.INIT = 1'b0;
  X_FF key1_45 (
    .I(key_45_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[45] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_46.INIT = 1'b0;
  X_FF key1_46 (
    .I(key_46_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[46] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_47.INIT = 1'b0;
  X_FF key1_47 (
    .I(key_47_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[47] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_48.INIT = 1'b0;
  X_FF key1_48 (
    .I(key_48_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[48] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd7_80.INIT = 1'b0;
  X_SFF state_FFd7_80 (
    .I(state_FFd8),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd7),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam key1_50.INIT = 1'b0;
  X_FF key1_50 (
    .I(key_50_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[50] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_51.INIT = 1'b0;
  X_FF key1_51 (
    .I(key_51_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[51] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_52.INIT = 1'b0;
  X_FF key1_52 (
    .I(key_52_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[52] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_53.INIT = 1'b0;
  X_FF key1_53 (
    .I(key_53_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[53] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_54.INIT = 1'b0;
  X_FF key1_54 (
    .I(key_54_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[54] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_55.INIT = 1'b0;
  X_FF key1_55 (
    .I(key_55_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[55] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_56.INIT = 1'b0;
  X_FF key1_56 (
    .I(key_56_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[56] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_58.INIT = 1'b0;
  X_FF key1_58 (
    .I(key_58_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[58] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_59.INIT = 1'b0;
  X_FF key1_59 (
    .I(key_59_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[59] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_60.INIT = 1'b0;
  X_FF key1_60 (
    .I(key_60_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[60] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_61.INIT = 1'b0;
  X_FF key1_61 (
    .I(key_61_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[61] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_62.INIT = 1'b0;
  X_FF key1_62 (
    .I(key_62_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[62] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam key1_63.INIT = 1'b0;
  X_FF key1_63 (
    .I(key_63_IBUF),
    .CE(_n0029),
    .CLK(clk_BUFGP),
    .O(\key1[63] ),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_1.INIT = 1'b0;
  X_FF data1_1 (
    .I(_n0013[0]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[1]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_2.INIT = 1'b0;
  X_FF data1_2 (
    .I(_n0013[1]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[2]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_3.INIT = 1'b0;
  X_FF data1_3 (
    .I(_n0013[2]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[3]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_4.INIT = 1'b0;
  X_FF data1_4 (
    .I(_n0013[3]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[4]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_5.INIT = 1'b0;
  X_FF data1_5 (
    .I(_n0013[4]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[5]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_6.INIT = 1'b0;
  X_FF data1_6 (
    .I(_n0013[5]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[6]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_7.INIT = 1'b0;
  X_FF data1_7 (
    .I(_n0013[6]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[7]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_8.INIT = 1'b0;
  X_FF data1_8 (
    .I(_n0013[7]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[8]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_9.INIT = 1'b0;
  X_FF data1_9 (
    .I(_n0013[8]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[9]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_10.INIT = 1'b0;
  X_FF data1_10 (
    .I(_n0013[9]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[10]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_11.INIT = 1'b0;
  X_FF data1_11 (
    .I(_n0013[10]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[11]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_12.INIT = 1'b0;
  X_FF data1_12 (
    .I(_n0013[11]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[12]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_13.INIT = 1'b0;
  X_FF data1_13 (
    .I(_n0013[12]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[13]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_14.INIT = 1'b0;
  X_FF data1_14 (
    .I(_n0013[13]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[14]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_15.INIT = 1'b0;
  X_FF data1_15 (
    .I(_n0013[14]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[15]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_16.INIT = 1'b0;
  X_FF data1_16 (
    .I(_n0013[15]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[16]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_17.INIT = 1'b0;
  X_FF data1_17 (
    .I(_n0013[16]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[17]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_18.INIT = 1'b0;
  X_FF data1_18 (
    .I(_n0013[17]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[18]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_19.INIT = 1'b0;
  X_FF data1_19 (
    .I(_n0013[18]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[19]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_20.INIT = 1'b0;
  X_FF data1_20 (
    .I(_n0013[19]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[20]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_21.INIT = 1'b0;
  X_FF data1_21 (
    .I(_n0013[20]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[21]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_22.INIT = 1'b0;
  X_FF data1_22 (
    .I(_n0013[21]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[22]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_23.INIT = 1'b0;
  X_FF data1_23 (
    .I(_n0013[22]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[23]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_24.INIT = 1'b0;
  X_FF data1_24 (
    .I(_n0013[23]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[24]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_25.INIT = 1'b0;
  X_FF data1_25 (
    .I(_n0013[24]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[25]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_26.INIT = 1'b0;
  X_FF data1_26 (
    .I(_n0013[25]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[26]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_27.INIT = 1'b0;
  X_FF data1_27 (
    .I(_n0013[26]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[27]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_28.INIT = 1'b0;
  X_FF data1_28 (
    .I(_n0013[27]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[28]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_29.INIT = 1'b0;
  X_FF data1_29 (
    .I(_n0013[28]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[29]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_30.INIT = 1'b0;
  X_FF data1_30 (
    .I(_n0013[29]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[30]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_31.INIT = 1'b0;
  X_FF data1_31 (
    .I(_n0013[30]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[31]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_32.INIT = 1'b0;
  X_FF data1_32 (
    .I(_n0013[31]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[32]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_33.INIT = 1'b0;
  X_FF data1_33 (
    .I(_n0013[32]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[33]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_34.INIT = 1'b0;
  X_FF data1_34 (
    .I(_n0013[33]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[34]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_35.INIT = 1'b0;
  X_FF data1_35 (
    .I(_n0013[34]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[35]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_36.INIT = 1'b0;
  X_FF data1_36 (
    .I(_n0013[35]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[36]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_37.INIT = 1'b0;
  X_FF data1_37 (
    .I(_n0013[36]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[37]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_38.INIT = 1'b0;
  X_FF data1_38 (
    .I(_n0013[37]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[38]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_39.INIT = 1'b0;
  X_FF data1_39 (
    .I(_n0013[38]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[39]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_40.INIT = 1'b0;
  X_FF data1_40 (
    .I(_n0013[39]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[40]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_41.INIT = 1'b0;
  X_FF data1_41 (
    .I(_n0013[40]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[41]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_42.INIT = 1'b0;
  X_FF data1_42 (
    .I(_n0013[41]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[42]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_43.INIT = 1'b0;
  X_FF data1_43 (
    .I(_n0013[42]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[43]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_44.INIT = 1'b0;
  X_FF data1_44 (
    .I(_n0013[43]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[44]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_45.INIT = 1'b0;
  X_FF data1_45 (
    .I(_n0013[44]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[45]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_46.INIT = 1'b0;
  X_FF data1_46 (
    .I(_n0013[45]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[46]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_47.INIT = 1'b0;
  X_FF data1_47 (
    .I(_n0013[46]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[47]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_48.INIT = 1'b0;
  X_FF data1_48 (
    .I(_n0013[47]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[48]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_49.INIT = 1'b0;
  X_FF data1_49 (
    .I(_n0013[48]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[49]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_50.INIT = 1'b0;
  X_FF data1_50 (
    .I(_n0013[49]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[50]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_51.INIT = 1'b0;
  X_FF data1_51 (
    .I(_n0013[50]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[51]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_52.INIT = 1'b0;
  X_FF data1_52 (
    .I(_n0013[51]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[52]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_53.INIT = 1'b0;
  X_FF data1_53 (
    .I(_n0013[52]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[53]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_54.INIT = 1'b0;
  X_FF data1_54 (
    .I(_n0013[53]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[54]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_55.INIT = 1'b0;
  X_FF data1_55 (
    .I(_n0013[54]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[55]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_56.INIT = 1'b0;
  X_FF data1_56 (
    .I(_n0013[55]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[56]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_57.INIT = 1'b0;
  X_FF data1_57 (
    .I(_n0013[56]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[57]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_58.INIT = 1'b0;
  X_FF data1_58 (
    .I(_n0013[57]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[58]),
    .SET(GND),
    .RST(GSR)
  );
  defparam data1_59.INIT = 1'b0;
  X_FF data1_59 (
    .I(_n0013[58]),
    .CE(rst_IBUF),
    .CLK(clk_BUFGP),
    .O(data1[59]),
    .SET(GND),
    .RST(GSR)
  );
  defparam state_FFd4_81.INIT = 1'b0;
  X_SFF state_FFd4_81 (
    .I(state_FFd6),
    .SRST(_n0032[2]),
    .CLK(clk_BUFGP),
    .O(state_FFd4),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  X_BUF datain_63_IBUF_82 (
    .I(datain[63]),
    .O(datain_63_IBUF)
  );
  defparam roundsel_4.INIT = 1'b1;
  X_SFF roundsel_4 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel[4]),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam \roundsel<1>_mmx_out851 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out851  (
    .ADR0(\key1[38] ),
    .ADR1(\key1[22] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out85 )
  );
  defparam \Maddsub__n0017_Mxor_Result<3>_Xo<0>1 .INIT = 16'h8001;
  X_LUT4 \Maddsub__n0017_Mxor_Result<3>_Xo<0>1  (
    .ADR0(state_FFd6),
    .ADR1(roundsel[1]),
    .ADR2(roundsel[2]),
    .ADR3(roundsel[3]),
    .O(\Maddsub__n0017_Mxor_Result<3>_Xo [0])
  );
  X_INV \_n0032<2>1_INV_0  (
    .I(rst_IBUF),
    .O(_n0032[2])
  );
  defparam \key2<28>12 .INIT = 16'hCA00;
  X_LUT4 \key2<28>12  (
    .ADR0(\key1[13] ),
    .ADR1(\key1[21] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_2_1),
    .O(CHOICE1823)
  );
  X_BUF datain_27_IBUF_83 (
    .I(datain[27]),
    .O(datain_27_IBUF)
  );
  X_BUF key_61_IBUF_84 (
    .I(key[61]),
    .O(key_61_IBUF)
  );
  X_BUF datain_29_IBUF_85 (
    .I(datain[29]),
    .O(datain_29_IBUF)
  );
  defparam \roundsel<1>_mmx_out871 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out871  (
    .ADR0(\key1[32] ),
    .ADR1(\key1[16] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out87 )
  );
  defparam \key2<9>133_SW0 .INIT = 16'h0075;
  X_LUT4 \key2<9>133_SW0  (
    .ADR0(roundsel_2_10),
    .ADR1(CHOICE1411),
    .ADR2(N5169),
    .ADR3(CHOICE1421),
    .O(N5093)
  );
  X_BUF flag_IBUF_86 (
    .I(flag),
    .O(flag_IBUF)
  );
  X_BUF datain_4_IBUF_87 (
    .I(datain[4]),
    .O(datain_4_IBUF)
  );
  defparam \roundsel<1>_mmx_out921 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out921  (
    .ADR0(\key1[24] ),
    .ADR1(\key1[16] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out92 )
  );
  X_BUF datain_31_IBUF_88 (
    .I(datain[31]),
    .O(datain_31_IBUF)
  );
  defparam \key2<15>133_SW0 .INIT = 16'h0705;
  X_LUT4 \key2<15>133_SW0  (
    .ADR0(roundsel_3_6),
    .ADR1(CHOICE585),
    .ADR2(CHOICE595),
    .ADR3(N5129),
    .O(N5095)
  );
  X_BUF datain_2_IBUF_89 (
    .I(datain[2]),
    .O(datain_2_IBUF)
  );
  X_BUF datain_22_IBUF_90 (
    .I(datain[22]),
    .O(datain_22_IBUF)
  );
  X_BUF datain_33_IBUF_91 (
    .I(datain[33]),
    .O(datain_33_IBUF)
  );
  X_BUF datain_35_IBUF_92 (
    .I(datain[35]),
    .O(datain_35_IBUF)
  );
  X_BUF datain_37_IBUF_93 (
    .I(datain[37]),
    .O(datain_37_IBUF)
  );
  defparam \key2<19>90 .INIT = 16'hFAF8;
  X_LUT4 \key2<19>90  (
    .ADR0(roundsel[4]),
    .ADR1(N5940),
    .ADR2(CHOICE867),
    .ADR3(CHOICE851),
    .O(\key2[19] )
  );
  X_BUF key_43_IBUF_94 (
    .I(key[43]),
    .O(key_43_IBUF)
  );
  defparam \roundsel<1>_mmx_out881 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out881  (
    .ADR0(\key1[48] ),
    .ADR1(\key1[64] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out88 )
  );
  defparam roundsel_4_2_95.INIT = 1'b1;
  X_SFF roundsel_4_2_95 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_2),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  X_BUF datain_39_IBUF_96 (
    .I(datain[39]),
    .O(datain_39_IBUF)
  );
  X_BUF datain_41_IBUF_97 (
    .I(datain[41]),
    .O(datain_41_IBUF)
  );
  X_BUF datain_6_IBUF_98 (
    .I(datain[6]),
    .O(datain_6_IBUF)
  );
  X_BUF datain_10_IBUF_99 (
    .I(datain[10]),
    .O(datain_10_IBUF)
  );
  defparam \key2<31>90 .INIT = 16'hFAF8;
  X_LUT4 \key2<31>90  (
    .ADR0(roundsel[4]),
    .ADR1(CHOICE1104),
    .ADR2(CHOICE1122),
    .ADR3(CHOICE1106),
    .O(\key2[31] )
  );
  X_BUF datain_60_IBUF_100 (
    .I(datain[60]),
    .O(datain_60_IBUF)
  );
  defparam \roundsel<1>_mmx_out931 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out931  (
    .ADR0(\key1[55] ),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out93 )
  );
  defparam \roundsel<1>_mmx_out911 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out911  (
    .ADR0(\key1[23] ),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out91 )
  );
  defparam \roundsel<1>_mmx_out891 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out891  (
    .ADR0(\key1[13] ),
    .ADR1(\key1[5] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out89 )
  );
  X_BUF datain_43_IBUF_101 (
    .I(datain[43]),
    .O(datain_43_IBUF)
  );
  defparam \roundsel<1>_mmx_out96 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out96  (
    .ADR0(\key1[8] ),
    .ADR1(\key1[21] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out9 )
  );
  X_BUF datain_45_IBUF_102 (
    .I(datain[45]),
    .O(datain_45_IBUF)
  );
  X_BUF datain_47_IBUF_103 (
    .I(datain[47]),
    .O(datain_47_IBUF)
  );
  defparam \roundsel<1>_mmx_out901 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out901  (
    .ADR0(\key1[16] ),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out90 )
  );
  defparam \key2<46>133_SW0 .INIT = 16'h0705;
  X_LUT4 \key2<46>133_SW0  (
    .ADR0(roundsel_2_13),
    .ADR1(CHOICE1887),
    .ADR2(CHOICE1897),
    .ADR3(N5139),
    .O(N5113)
  );
  defparam \roundsel<1>_mmx_out951 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out951  (
    .ADR0(\key1[30] ),
    .ADR1(\key1[46] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out95 )
  );
  defparam roundsel_3_16_104.INIT = 1'b1;
  X_SFF roundsel_3_16_104 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_16),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam \key2<17>133_SW0 .INIT = 16'h005D;
  X_LUT4 \key2<17>133_SW0  (
    .ADR0(roundsel_3_6),
    .ADR1(N5141),
    .ADR2(CHOICE521),
    .ADR3(CHOICE531),
    .O(N5097)
  );
  defparam \roundsel<1>_mmx_out2 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out2  (
    .ADR0(\key1[13] ),
    .ADR1(\key1[62] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out )
  );
  defparam \roundsel<1>_mmx_out12 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out12  (
    .ADR0(\key1[8] ),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out1 )
  );
  defparam \roundsel<1>_mmx_out101 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out101  (
    .ADR0(\key1[31] ),
    .ADR1(\key1[15] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out10 )
  );
  defparam \roundsel<1>_mmx_out111 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out111  (
    .ADR0(\key1[47] ),
    .ADR1(\key1[55] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out11 )
  );
  defparam \roundsel<1>_mmx_out121 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out121  (
    .ADR0(\key1[64] ),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out12 )
  );
  defparam \roundsel<1>_mmx_out131 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out131  (
    .ADR0(\key1[63] ),
    .ADR1(\key1[47] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out13 )
  );
  defparam \roundsel<1>_mmx_out141 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out141  (
    .ADR0(\key1[40] ),
    .ADR1(\key1[48] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out14 )
  );
  defparam \roundsel<1>_mmx_out151 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out151  (
    .ADR0(\key1[14] ),
    .ADR1(\key1[30] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out15 )
  );
  defparam \roundsel<1>_mmx_out161 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out161  (
    .ADR0(\key1[54] ),
    .ADR1(\key1[46] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out16 )
  );
  defparam \roundsel<1>_mmx_out171 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out171  (
    .ADR0(\key1[30] ),
    .ADR1(\key1[38] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out17 )
  );
  defparam \roundsel<1>_mmx_out181 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out181  (
    .ADR0(\key1[31] ),
    .ADR1(\key1[23] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out18 )
  );
  defparam \roundsel<1>_mmx_out191 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out191  (
    .ADR0(\key1[15] ),
    .ADR1(\key1[7] ),
    .ADR2(roundsel_1_6),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out19 )
  );
  defparam \roundsel<1>_mmx_out22 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out22  (
    .ADR0(\key1[48] ),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out2 )
  );
  defparam \roundsel<1>_mmx_out201 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out201  (
    .ADR0(\key1[24] ),
    .ADR1(\key1[40] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out20 )
  );
  defparam \roundsel<1>_mmx_out211 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out211  (
    .ADR0(\key1[62] ),
    .ADR1(\key1[46] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out21 )
  );
  defparam \roundsel<1>_mmx_out221 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out221  (
    .ADR0(\key1[24] ),
    .ADR1(\key1[32] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out22 )
  );
  defparam \roundsel<1>_mmx_out231 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out231  (
    .ADR0(\key1[13] ),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out23 )
  );
  defparam \roundsel<1>_mmx_out241 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out241  (
    .ADR0(\key1[20] ),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out24 )
  );
  defparam \roundsel<1>_mmx_out251 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out251  (
    .ADR0(\key1[52] ),
    .ADR1(\key1[36] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out25 )
  );
  defparam \roundsel<1>_mmx_out261 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out261  (
    .ADR0(\key1[37] ),
    .ADR1(\key1[53] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out26 )
  );
  defparam \roundsel<1>_mmx_out271 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out271  (
    .ADR0(\key1[10] ),
    .ADR1(\key1[61] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out27 )
  );
  defparam \roundsel<1>_mmx_out281 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out281  (
    .ADR0(\key1[42] ),
    .ADR1(\key1[26] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out28 )
  );
  defparam \roundsel<1>_mmx_out291 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out291  (
    .ADR0(\key1[58] ),
    .ADR1(\key1[11] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out29 )
  );
  defparam \roundsel<1>_mmx_out32 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out32  (
    .ADR0(\key1[22] ),
    .ADR1(\key1[6] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out3 )
  );
  defparam \roundsel<1>_mmx_out301 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out301  (
    .ADR0(\key1[35] ),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_1_6),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out30 )
  );
  defparam \roundsel<1>_mmx_out311 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out311  (
    .ADR0(\key1[24] ),
    .ADR1(\key1[8] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out31 )
  );
  defparam \roundsel<1>_mmx_out321 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out321  (
    .ADR0(\key1[35] ),
    .ADR1(\key1[19] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out32 )
  );
  defparam \roundsel<1>_mmx_out331 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out331  (
    .ADR0(\key1[51] ),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out33 )
  );
  defparam \roundsel<1>_mmx_out341 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out341  (
    .ADR0(\key1[20] ),
    .ADR1(\key1[36] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out34 )
  );
  defparam \roundsel<1>_mmx_out351 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out351  (
    .ADR0(\key1[60] ),
    .ADR1(\key1[52] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out35 )
  );
  defparam \roundsel<1>_mmx_out361 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out361  (
    .ADR0(\key1[34] ),
    .ADR1(\key1[26] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out36 )
  );
  defparam \roundsel<1>_mmx_out371 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out371  (
    .ADR0(\key1[3] ),
    .ADR1(\key1[50] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out37 )
  );
  defparam \roundsel<1>_mmx_out381 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out381  (
    .ADR0(\key1[28] ),
    .ADR1(\key1[12] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out38 )
  );
  defparam \roundsel<1>_mmx_out391 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out391  (
    .ADR0(\key1[60] ),
    .ADR1(\key1[44] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out39 )
  );
  defparam \roundsel<1>_mmx_out410 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out410  (
    .ADR0(\key1[40] ),
    .ADR1(\key1[32] ),
    .ADR2(roundsel_1_14),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out4 )
  );
  defparam \roundsel<1>_mmx_out401 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out401  (
    .ADR0(\key1[40] ),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out40 )
  );
  defparam \roundsel<1>_mmx_out411 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out411  (
    .ADR0(\key1[61] ),
    .ADR1(\key1[45] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out41 )
  );
  defparam \roundsel<1>_mmx_out421 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out421  (
    .ADR0(\key1[10] ),
    .ADR1(\key1[18] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out42 )
  );
  defparam \roundsel<1>_mmx_out431 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out431  (
    .ADR0(\key1[19] ),
    .ADR1(\key1[11] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out43 )
  );
  defparam \roundsel<1>_mmx_out441 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out441  (
    .ADR0(\key1[35] ),
    .ADR1(\key1[51] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out44 )
  );
  defparam \roundsel<1>_mmx_out451 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out451  (
    .ADR0(\key1[45] ),
    .ADR1(\key1[60] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out45 )
  );
  defparam \roundsel<1>_mmx_out461 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out461  (
    .ADR0(\key1[28] ),
    .ADR1(\key1[36] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out46 )
  );
  defparam \roundsel<1>_mmx_out471 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out471  (
    .ADR0(\key1[37] ),
    .ADR1(\key1[52] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out47 )
  );
  defparam \roundsel<1>_mmx_out481 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out481  (
    .ADR0(\key1[53] ),
    .ADR1(\key1[2] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out48 )
  );
  defparam \roundsel<1>_mmx_out491 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out491  (
    .ADR0(\key1[34] ),
    .ADR1(\key1[18] ),
    .ADR2(roundsel_11),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out49 )
  );
  defparam \roundsel<1>_mmx_out52 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out52  (
    .ADR0(\key1[7] ),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out5 )
  );
  defparam \roundsel<1>_mmx_out501 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out501  (
    .ADR0(\key1[58] ),
    .ADR1(\key1[42] ),
    .ADR2(roundsel_1_4),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out50 )
  );
  defparam \roundsel<1>_mmx_out511 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out511  (
    .ADR0(\key1[27] ),
    .ADR1(\key1[11] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out51 )
  );
  defparam \roundsel<1>_mmx_out531 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out531  (
    .ADR0(\key1[12] ),
    .ADR1(\key1[20] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out53 )
  );
  defparam \roundsel<1>_mmx_out541 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out541  (
    .ADR0(\key1[61] ),
    .ADR1(\key1[2] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out54 )
  );
  defparam \roundsel<1>_mmx_out551 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out551  (
    .ADR0(\key1[23] ),
    .ADR1(\key1[7] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out55 )
  );
  defparam \roundsel<1>_mmx_out561 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out561  (
    .ADR0(\key1[45] ),
    .ADR1(\key1[53] ),
    .ADR2(roundsel_12),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out56 )
  );
  defparam \roundsel<1>_mmx_out581 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out581  (
    .ADR0(\key1[10] ),
    .ADR1(\key1[2] ),
    .ADR2(roundsel_1_22),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out58 )
  );
  defparam \roundsel<1>_mmx_out591 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out591  (
    .ADR0(\key1[35] ),
    .ADR1(\key1[43] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out59 )
  );
  defparam \roundsel<1>_mmx_out610 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out610  (
    .ADR0(\key1[63] ),
    .ADR1(\key1[55] ),
    .ADR2(roundsel_1_14),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out6 )
  );
  defparam \roundsel<1>_mmx_out601 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out601  (
    .ADR0(\key1[59] ),
    .ADR1(\key1[12] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out60 )
  );
  defparam \roundsel<1>_mmx_out611 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out611  (
    .ADR0(\key1[44] ),
    .ADR1(\key1[28] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out61 )
  );
  defparam \roundsel<1>_mmx_out641 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out641  (
    .ADR0(\key1[47] ),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out64 )
  );
  defparam \roundsel<1>_mmx_out651 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out651  (
    .ADR0(\key1[18] ),
    .ADR1(\key1[2] ),
    .ADR2(roundsel_1_19),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out65 )
  );
  defparam \roundsel<1>_mmx_out661 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out661  (
    .ADR0(\key1[43] ),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out66 )
  );
  defparam \roundsel<1>_mmx_out671 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out671  (
    .ADR0(\key1[19] ),
    .ADR1(\key1[3] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out67 )
  );
  defparam \roundsel<1>_mmx_out681 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out681  (
    .ADR0(\key1[44] ),
    .ADR1(\key1[36] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out68 )
  );
  defparam \roundsel<1>_mmx_out691 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out691  (
    .ADR0(\key1[28] ),
    .ADR1(\key1[20] ),
    .ADR2(roundsel_1_14),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out69 )
  );
  defparam \roundsel<1>_mmx_out71 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out71  (
    .ADR0(\key1[8] ),
    .ADR1(\key1[16] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out7 )
  );
  defparam \roundsel<1>_mmx_out701 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out701  (
    .ADR0(\key1[12] ),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_1_14),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out70 )
  );
  defparam \roundsel<1>_mmx_out711 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out711  (
    .ADR0(\key1[59] ),
    .ADR1(\key1[51] ),
    .ADR2(roundsel_1_15),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out71 )
  );
  defparam \roundsel<1>_mmx_out721 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out721  (
    .ADR0(\key1[34] ),
    .ADR1(\key1[50] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out72 )
  );
  defparam \roundsel<1>_mmx_out731 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out731  (
    .ADR0(\key1[10] ),
    .ADR1(\key1[26] ),
    .ADR2(roundsel_11),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out73 )
  );
  defparam \roundsel<1>_mmx_out741 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out741  (
    .ADR0(\key1[58] ),
    .ADR1(\key1[50] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out74 )
  );
  defparam \roundsel<1>_mmx_out761 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out761  (
    .ADR0(\key1[14] ),
    .ADR1(\key1[22] ),
    .ADR2(roundsel_1_21),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out76 )
  );
  defparam \roundsel<1>_mmx_out771 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out771  (
    .ADR0(\key1[54] ),
    .ADR1(\key1[38] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out77 )
  );
  defparam \roundsel<1>_mmx_out781 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out781  (
    .ADR0(\key1[21] ),
    .ADR1(\key1[5] ),
    .ADR2(roundsel_1_16),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out78 )
  );
  defparam \roundsel<1>_mmx_out791 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out791  (
    .ADR0(\key1[48] ),
    .ADR1(\key1[32] ),
    .ADR2(roundsel_1_17),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out79 )
  );
  defparam \roundsel<1>_mmx_out801 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out801  (
    .ADR0(\key1[15] ),
    .ADR1(\key1[64] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out80 )
  );
  defparam \roundsel<1>_mmx_out811 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out811  (
    .ADR0(\key1[47] ),
    .ADR1(\key1[31] ),
    .ADR2(roundsel_1_20),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out81 )
  );
  defparam \roundsel<1>_mmx_out821 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out821  (
    .ADR0(\key1[63] ),
    .ADR1(\key1[6] ),
    .ADR2(roundsel_1_8),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out82 )
  );
  defparam \roundsel<1>_mmx_out831 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out831  (
    .ADR0(\key1[31] ),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_1_18),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out83 )
  );
  X_BUF key_39_IBUF_105 (
    .I(key[39]),
    .O(key_39_IBUF)
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_23 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_23  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_46 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_47 ),
    .O(\c1/u5/Mrom_dout_N10 )
  );
  X_BUF dataout_46_OBUF (
    .I(dataout_46),
    .O(\dataout_46_OBUF.GTS.TRI )
  );
  X_BUF dataout_27_OBUF (
    .I(dataout_27),
    .O(\dataout_27_OBUF.GTS.TRI )
  );
  X_BUF dataout_34_OBUF (
    .I(dataout_34),
    .O(\dataout_34_OBUF.GTS.TRI )
  );
  X_BUF dataout_50_OBUF (
    .I(dataout_50),
    .O(\dataout_50_OBUF.GTS.TRI )
  );
  X_BUF dataout_33_OBUF (
    .I(dataout_33),
    .O(\dataout_33_OBUF.GTS.TRI )
  );
  X_BUF dataout_40_OBUF (
    .I(dataout_40),
    .O(\dataout_40_OBUF.GTS.TRI )
  );
  X_BUF dataout_44_OBUF (
    .I(dataout_44),
    .O(\dataout_44_OBUF.GTS.TRI )
  );
  X_BUF dataout_24_OBUF (
    .I(dataout_24),
    .O(\dataout_24_OBUF.GTS.TRI )
  );
  defparam \c1/Mxor_OUTR_Result<3>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<3>1  (
    .ADR0(\c1/X[36] ),
    .ADR1(data1[36]),
    .ADR2(\c1/u5/Mrom_dout_N3 ),
    .ADR3(\c1/u5/Mrom_dout_N4 ),
    .O(cipherout2[4])
  );
  defparam \_n0013<14>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<14>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[53]),
    .ADR2(state_FFd8),
    .ADR3(datain_15_IBUF),
    .O(CHOICE1038)
  );
  X_BUF dataout_9_OBUF (
    .I(dataout_9),
    .O(\dataout_9_OBUF.GTS.TRI )
  );
  X_BUF datain_38_IBUF_106 (
    .I(datain[38]),
    .O(datain_38_IBUF)
  );
  X_BUF key_7_IBUF_107 (
    .I(key[7]),
    .O(key_7_IBUF)
  );
  defparam \c1/Mxor_OUTR_Result<19>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<19>1  (
    .ADR0(\c1/X[12] ),
    .ADR1(data1[52]),
    .ADR2(\c1/u1/Mrom_dout_N0 ),
    .ADR3(\c1/u1/Mrom_dout_N1 ),
    .O(cipherout2[20])
  );
  defparam \_n0013<11>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<11>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[29]),
    .ADR2(state_FFd8),
    .ADR3(datain_12_IBUF),
    .O(CHOICE1936)
  );
  X_BUF key_59_IBUF_108 (
    .I(key[59]),
    .O(key_59_IBUF)
  );
  X_BUF key_35_IBUF_109 (
    .I(key[35]),
    .O(key_35_IBUF)
  );
  defparam \c1/Mxor_OUTR_Result<31>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<31>1  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[64]),
    .ADR2(\c1/u3/Mrom_dout_N9 ),
    .ADR3(\c1/u3/Mrom_dout_N10 ),
    .O(cipherout2[32])
  );
  defparam \_n0013<11>6 .INIT = 4'h8;
  X_LUT2 \_n0013<11>6  (
    .ADR0(data1[12]),
    .ADR1(N01),
    .O(CHOICE1937)
  );
  X_BUF key_28_IBUF_110 (
    .I(key[28]),
    .O(key_28_IBUF)
  );
  defparam \c1/Mxor_X_Result<5>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<5>1  (
    .ADR0(data1[28]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE339),
    .ADR3(N5153),
    .O(\c1/X[6] )
  );
  X_BUF datain_57_IBUF_111 (
    .I(datain[57]),
    .O(datain_57_IBUF)
  );
  X_BUF datain_59_IBUF_112 (
    .I(datain[59]),
    .O(datain_59_IBUF)
  );
  defparam \c1/Mxor_X_Result<11>1 .INIT = 16'h6636;
  X_LUT4 \c1/Mxor_X_Result<11>1  (
    .ADR0(CHOICE283),
    .ADR1(data1[24]),
    .ADR2(roundsel[4]),
    .ADR3(N5171),
    .O(\c1/X[12] )
  );
  defparam \c1/Mxor_X_Result<12>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<12>1  (
    .ADR0(data1[25]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE491),
    .ADR3(N5115),
    .O(\c1/X[13] )
  );
  X_BUF datain_3_IBUF_113 (
    .I(datain[3]),
    .O(datain_3_IBUF)
  );
  defparam \c1/Mxor_X_Result<17>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<17>1  (
    .ADR0(data1[20]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE259),
    .ADR3(N5179),
    .O(\c1/X[18] )
  );
  defparam \c1/Mxor_X_Result<18>1 .INIT = 16'h6636;
  X_LUT4 \c1/Mxor_X_Result<18>1  (
    .ADR0(CHOICE867),
    .ADR1(data1[21]),
    .ADR2(roundsel[4]),
    .ADR3(N5181),
    .O(\c1/X[19] )
  );
  defparam \c1/Mxor_X_Result<20>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<20>1  (
    .ADR0(data1[19]),
    .ADR1(roundsel[3]),
    .ADR2(CHOICE996),
    .ADR3(N5099),
    .O(\c1/X[21] )
  );
  defparam \c1/Mxor_X_Result<23>1 .INIT = 16'h6636;
  X_LUT4 \c1/Mxor_X_Result<23>1  (
    .ADR0(CHOICE431),
    .ADR1(data1[16]),
    .ADR2(roundsel[4]),
    .ADR3(N5123),
    .O(\c1/X[24] )
  );
  defparam \c1/Mxor_X_Result<24>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<24>1  (
    .ADR0(data1[17]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1150),
    .ADR3(N5117),
    .O(\c1/X[25] )
  );
  X_BUF datain_5_IBUF_114 (
    .I(datain[5]),
    .O(datain_5_IBUF)
  );
  defparam \c1/Mxor_X_Result<26>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<26>1  (
    .ADR0(data1[15]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1340),
    .ADR3(N5101),
    .O(\c1/X[27] )
  );
  defparam \c1/Mxor_X_Result<27>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<27>1  (
    .ADR0(data1[14]),
    .ADR1(roundsel[3]),
    .ADR2(CHOICE1849),
    .ADR3(N5103),
    .O(\c1/X[28] )
  );
  defparam \c1/Mxor_X_Result<29>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<29>1  (
    .ADR0(data1[12]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE463),
    .ADR3(N5155),
    .O(\c1/X[30] )
  );
  X_BUF datain_56_IBUF_115 (
    .I(datain[56]),
    .O(datain_56_IBUF)
  );
  X_BUF datain_61_IBUF_116 (
    .I(datain[61]),
    .O(datain_61_IBUF)
  );
  defparam \c1/Mxor_X_Result<35>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<35>1  (
    .ADR0(data1[8]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE399),
    .ADR3(N5157),
    .O(\c1/X[36] )
  );
  defparam \c1/Mxor_X_Result<36>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<36>1  (
    .ADR0(data1[9]),
    .ADR1(roundsel[4]),
    .ADR2(N5119),
    .ADR3(CHOICE1178),
    .O(\c1/X[37] )
  );
  defparam \c1/Mxor_X_Result<41>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<41>1  (
    .ADR0(data1[4]),
    .ADR1(roundsel[4]),
    .ADR2(N5125),
    .ADR3(CHOICE311),
    .O(\c1/X[42] )
  );
  defparam \c1/Mxor_X_Result<42>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<42>1  (
    .ADR0(data1[5]),
    .ADR1(roundsel[4]),
    .ADR2(N5121),
    .ADR3(CHOICE1206),
    .O(\c1/X[43] )
  );
  defparam \c1/Mxor_X_Result<44>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<44>1  (
    .ADR0(data1[3]),
    .ADR1(roundsel[3]),
    .ADR2(CHOICE1881),
    .ADR3(N5111),
    .O(\c1/X[45] )
  );
  defparam \c1/Mxor_X_Result<47>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<47>1  (
    .ADR0(data1[32]),
    .ADR1(roundsel[4]),
    .ADR2(N5159),
    .ADR3(CHOICE367),
    .O(\c1/X[48] )
  );
  X_BUF datain_7_IBUF_117 (
    .I(datain[7]),
    .O(datain_7_IBUF)
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_01 .INIT = 16'h9E61;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_01  (
    .ADR0(\c1/X[45] ),
    .ADR1(\c1/X[44] ),
    .ADR2(\c1/X[47] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_0 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_16 .INIT = 16'h529B;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_16  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[45] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_1 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_21 .INIT = 16'h4DA3;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_21  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[45] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_2 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_31 .INIT = 16'hA6C6;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_31  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[46] ),
    .ADR3(\c1/X[45] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_3 )
  );
  X_BUF dataout_47_OBUF (
    .I(dataout_47),
    .O(\dataout_47_OBUF.GTS.TRI )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_41 .INIT = 16'h9C36;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_41  (
    .ADR0(N5933),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[46] ),
    .ADR3(\c1/X[45] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_4 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_51 .INIT = 16'hD398;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_51  (
    .ADR0(\c1/X[45] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[44] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_5 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_61 .INIT = 16'h6659;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_61  (
    .ADR0(\c1/X[45] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[44] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_6 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_71 .INIT = 16'hC635;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_71  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[45] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_7 )
  );
  X_BUF dataout_41_OBUF (
    .I(dataout_41),
    .O(\dataout_41_OBUF.GTS.TRI )
  );
  defparam \c1/Mxor_OUTR_Result<17>1_F_SW0 .INIT = 16'h652E;
  X_LUT4 \c1/Mxor_OUTR_Result<17>1_F_SW0  (
    .ADR0(\c1/X[45] ),
    .ADR1(\c1/X[47] ),
    .ADR2(N5934),
    .ADR3(\c1/X[44] ),
    .O(N5490)
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_101 .INIT = 16'h1EA5;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_101  (
    .ADR0(N5935),
    .ADR1(\c1/X[45] ),
    .ADR2(\c1/X[44] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_10 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_111 .INIT = 16'h693C;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_111  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[45] ),
    .ADR2(\c1/X[47] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_11 )
  );
  X_BUF dataout_45_OBUF (
    .I(dataout_45),
    .O(\dataout_45_OBUF.GTS.TRI )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_121 .INIT = 16'h4B65;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_121  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[45] ),
    .ADR2(\c1/X[46] ),
    .ADR3(\c1/X[47] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_12 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_131 .INIT = 16'h49B6;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_131  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[47] ),
    .ADR2(\c1/X[45] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_13 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_141 .INIT = 16'h9C72;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_141  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[45] ),
    .ADR2(\c1/X[46] ),
    .ADR3(\c1/X[47] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_14 )
  );
  defparam \c1/u7/Mrom_dout_inst_lut4_151 .INIT = 16'h8E74;
  X_LUT4 \c1/u7/Mrom_dout_inst_lut4_151  (
    .ADR0(\c1/X[44] ),
    .ADR1(\c1/X[45] ),
    .ADR2(\c1/X[47] ),
    .ADR3(\c1/X[46] ),
    .O(\c1/u7/Mrom_dout_inst_lut4_15 )
  );
  X_BUF dataout_43_OBUF (
    .I(dataout_43),
    .O(\dataout_43_OBUF.GTS.TRI )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_62 .INIT = 16'h64B9;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_62  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(N5187),
    .ADR3(N5186),
    .O(\c1/u1/Mrom_dout_N9 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_161 .INIT = 16'h9D92;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_161  (
    .ADR0(\c1/X[38] ),
    .ADR1(\c1/X[39] ),
    .ADR2(\c1/X[40] ),
    .ADR3(\c1/X[41] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_16 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_171 .INIT = 16'h526B;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_171  (
    .ADR0(\c1/X[39] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[38] ),
    .ADR3(\c1/X[41] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_17 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_181 .INIT = 16'h586B;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_181  (
    .ADR0(\c1/X[39] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[38] ),
    .ADR3(\c1/X[41] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_18 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_191 .INIT = 16'h6396;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_191  (
    .ADR0(\c1/X[41] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[39] ),
    .ADR3(\c1/X[38] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_19 )
  );
  X_BUF dataout_51_OBUF (
    .I(dataout_51),
    .O(\dataout_51_OBUF.GTS.TRI )
  );
  X_BUF key_64_IBUF_118 (
    .I(key[64]),
    .O(key_64_IBUF)
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_241 .INIT = 16'h6A59;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_241  (
    .ADR0(N5929),
    .ADR1(\c1/X[41] ),
    .ADR2(\c1/X[40] ),
    .ADR3(\c1/X[39] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_24 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_251 .INIT = 16'hB295;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_251  (
    .ADR0(\c1/X[38] ),
    .ADR1(\c1/X[40] ),
    .ADR2(N5932),
    .ADR3(\c1/X[39] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_25 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_261 .INIT = 16'h3D62;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_261  (
    .ADR0(N5931),
    .ADR1(\c1/X[41] ),
    .ADR2(\c1/X[39] ),
    .ADR3(\c1/X[38] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_26 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_271 .INIT = 16'hA969;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_271  (
    .ADR0(\c1/X[38] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[39] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_27 )
  );
  X_BUF key_45_IBUF_119 (
    .I(key[45]),
    .O(key_45_IBUF)
  );
  X_BUF dataout_42_OBUF (
    .I(dataout_42),
    .O(\dataout_42_OBUF.GTS.TRI )
  );
  X_BUF dataout_2_OBUF (
    .I(dataout_2),
    .O(\dataout_2_OBUF.GTS.TRI )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_291 .INIT = 16'h6999;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_291  (
    .ADR0(\c1/X[38] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[39] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_29 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_301 .INIT = 16'h49BC;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_301  (
    .ADR0(\c1/X[38] ),
    .ADR1(N5930),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[40] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_30 )
  );
  defparam \c1/u6/Mrom_dout_inst_lut4_311 .INIT = 16'h949E;
  X_LUT4 \c1/u6/Mrom_dout_inst_lut4_311  (
    .ADR0(\c1/X[38] ),
    .ADR1(\c1/X[39] ),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[40] ),
    .O(\c1/u6/Mrom_dout_inst_lut4_31 )
  );
  defparam \key2<28>25_SW0 .INIT = 16'hFF53;
  X_LUT4 \key2<28>25_SW0  (
    .ADR0(\key1[62] ),
    .ADR1(\key1[46] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_22),
    .O(N5135)
  );
  X_BUF key_52_IBUF_120 (
    .I(key[52]),
    .O(key_52_IBUF)
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_331 .INIT = 16'h6D62;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_331  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_33 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_351 .INIT = 16'h9C36;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_351  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[35] ),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[33] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_35 )
  );
  defparam \c1/u3/Mrom_dout_inst_mux_f5_39 .INIT = 16'hF690;
  X_LUT4 \c1/u3/Mrom_dout_inst_mux_f5_39  (
    .ADR0(data1[21]),
    .ADR1(\key2[19] ),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_78 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_74 ),
    .O(\c1/u3/Mrom_dout_N10 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_16 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_16  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_32 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_33 ),
    .O(\c1/u5/Mrom_dout_N0 )
  );
  X_BUF dataout_48_OBUF (
    .I(dataout_48),
    .O(\dataout_48_OBUF.GTS.TRI )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_361 .INIT = 16'hB64C;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_361  (
    .ADR0(\c1/X[32] ),
    .ADR1(N5926),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_36 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_371 .INIT = 16'h619B;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_371  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(N5927),
    .O(\c1/u5/Mrom_dout_inst_lut4_37 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_391 .INIT = 16'h2D66;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_391  (
    .ADR0(\c1/X[33] ),
    .ADR1(N5928),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[32] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_39 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_17 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_17  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_34 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_35 ),
    .O(\c1/u5/Mrom_dout_N1 )
  );
  X_BUF dataout_36_OBUF (
    .I(dataout_36),
    .O(\dataout_36_OBUF.GTS.TRI )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_411 .INIT = 16'h2D36;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_411  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[35] ),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[33] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_41 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_431 .INIT = 16'h96C9;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_431  (
    .ADR0(\c1/X[33] ),
    .ADR1(\c1/X[32] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_43 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_19 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_19  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_38 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_39 ),
    .O(\c1/u5/Mrom_dout_N4 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_20 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_20  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_40 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_41 ),
    .O(\c1/u5/Mrom_dout_N6 )
  );
  X_BUF dataout_31_OBUF (
    .I(dataout_31),
    .O(\dataout_31_OBUF.GTS.TRI )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_451 .INIT = 16'hA6C3;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_451  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_45 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_471 .INIT = 16'hCD38;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_471  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_47 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_21 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_21  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_42 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_43 ),
    .O(\c1/u5/Mrom_dout_N7 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_22 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_22  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_44 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_45 ),
    .O(\c1/u5/Mrom_dout_N9 )
  );
  X_BUF dataout_32_OBUF (
    .I(dataout_32),
    .O(\dataout_32_OBUF.GTS.TRI )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_521 .INIT = 16'h73C1;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_521  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[29] ),
    .ADR2(\c1/X[27] ),
    .ADR3(\c1/X[28] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_52 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_531 .INIT = 16'h86D3;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_531  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[29] ),
    .ADR2(\c1/X[27] ),
    .ADR3(\c1/X[28] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_53 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_541 .INIT = 16'h949E;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_541  (
    .ADR0(\c1/X[29] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[26] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_54 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_551 .INIT = 16'h946B;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_551  (
    .ADR0(\c1/X[29] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[26] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_55 )
  );
  defparam \_n0013<3>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<3>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[31]),
    .ADR2(state_FFd8),
    .ADR3(datain_4_IBUF),
    .O(CHOICE1345)
  );
  X_BUF dataout_29_OBUF (
    .I(dataout_29),
    .O(\dataout_29_OBUF.GTS.TRI )
  );
  X_BUF dataout_25_OBUF (
    .I(dataout_25),
    .O(\dataout_25_OBUF.GTS.TRI )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_601 .INIT = 16'hAC5A;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_601  (
    .ADR0(N5925),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[26] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_60 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_611 .INIT = 16'h7863;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_611  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[27] ),
    .ADR3(\c1/X[29] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_61 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_621 .INIT = 16'hA36C;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_621  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[29] ),
    .ADR2(\c1/X[27] ),
    .ADR3(\c1/X[28] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_62 )
  );
  defparam \c1/u4/Mrom_dout_inst_lut4_631 .INIT = 16'h296B;
  X_LUT4 \c1/u4/Mrom_dout_inst_lut4_631  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[29] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_lut4_63 )
  );
  X_BUF dataout_17_OBUF (
    .I(dataout_17),
    .O(\dataout_17_OBUF.GTS.TRI )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_641 .INIT = 16'hB41B;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_641  (
    .ADR0(\c1/X[23] ),
    .ADR1(\c1/X[22] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_64 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_651 .INIT = 16'hB169;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_651  (
    .ADR0(\c1/X[22] ),
    .ADR1(\c1/X[23] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_65 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_661 .INIT = 16'h267C;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_661  (
    .ADR0(\c1/X[22] ),
    .ADR1(\c1/X[23] ),
    .ADR2(\c1/X[21] ),
    .ADR3(\c1/X[20] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_66 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_671 .INIT = 16'h26D3;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_671  (
    .ADR0(\c1/X[23] ),
    .ADR1(\c1/X[22] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_67 )
  );
  defparam \key2<9>25_SW0 .INIT = 16'hF5F3;
  X_LUT4 \key2<9>25_SW0  (
    .ADR0(\key1[36] ),
    .ADR1(\key1[20] ),
    .ADR2(roundsel_3_5),
    .ADR3(roundsel_1_6),
    .O(N5169)
  );
  X_BUF key_62_IBUF_121 (
    .I(key[62]),
    .O(key_62_IBUF)
  );
  X_BUF dataout_3_OBUF (
    .I(dataout_3),
    .O(\dataout_3_OBUF.GTS.TRI )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_691 .INIT = 16'h2DE2;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_691  (
    .ADR0(\c1/X[22] ),
    .ADR1(\c1/X[23] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_69 )
  );
  X_BUF dataout_4_OBUF (
    .I(dataout_4),
    .O(\dataout_4_OBUF.GTS.TRI )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_711 .INIT = 16'hC9A3;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_711  (
    .ADR0(\c1/X[20] ),
    .ADR1(\c1/X[23] ),
    .ADR2(\c1/X[21] ),
    .ADR3(\c1/X[22] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_71 )
  );
  X_BUF key_63_IBUF_122 (
    .I(key[63]),
    .O(key_63_IBUF)
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_721 .INIT = 16'hC9A3;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_721  (
    .ADR0(N5922),
    .ADR1(\c1/X[23] ),
    .ADR2(\c1/X[22] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_72 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_731 .INIT = 16'h3867;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_731  (
    .ADR0(\c1/X[23] ),
    .ADR1(\c1/X[22] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_73 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_741 .INIT = 16'hE41E;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_741  (
    .ADR0(\c1/X[23] ),
    .ADR1(N5923),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_74 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_751 .INIT = 16'h96B8;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_751  (
    .ADR0(\c1/X[23] ),
    .ADR1(\c1/X[22] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_75 )
  );
  X_BUF datain_12_IBUF_123 (
    .I(datain[12]),
    .O(datain_12_IBUF)
  );
  X_BUF datain_1_IBUF_124 (
    .I(datain[1]),
    .O(datain_1_IBUF)
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_761 .INIT = 16'hC798;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_761  (
    .ADR0(N5924),
    .ADR1(\c1/X[22] ),
    .ADR2(\c1/X[20] ),
    .ADR3(\c1/X[21] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_76 )
  );
  X_BUF dataout_5_OBUF (
    .I(dataout_5),
    .O(\dataout_5_OBUF.GTS.TRI )
  );
  X_BUF dataout_6_OBUF (
    .I(dataout_6),
    .O(\dataout_6_OBUF.GTS.TRI )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_801 .INIT = 16'h5A3C;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_801  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_80 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_811 .INIT = 16'hA5C3;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_811  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_81 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_821 .INIT = 16'h9639;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_821  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_82 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_831 .INIT = 16'h7A25;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_831  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_83 )
  );
  X_BUF dataout_26_OBUF (
    .I(dataout_26),
    .O(\dataout_26_OBUF.GTS.TRI )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_841 .INIT = 16'h5A2B;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_841  (
    .ADR0(\c1/X[16] ),
    .ADR1(N5921),
    .ADR2(\c1/X[14] ),
    .ADR3(\c1/X[15] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_84 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_851 .INIT = 16'h69A6;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_851  (
    .ADR0(\c1/X[16] ),
    .ADR1(N5919),
    .ADR2(\c1/X[15] ),
    .ADR3(\c1/X[17] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_85 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_861 .INIT = 16'hA3D8;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_861  (
    .ADR0(\c1/X[16] ),
    .ADR1(N5920),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_86 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_871 .INIT = 16'h6C5A;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_871  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[17] ),
    .ADR2(\c1/X[14] ),
    .ADR3(\c1/X[15] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_87 )
  );
  X_BUF dataout_53_OBUF (
    .I(dataout_53),
    .O(\dataout_53_OBUF.GTS.TRI )
  );
  X_BUF dataout_28_OBUF (
    .I(dataout_28),
    .O(\dataout_28_OBUF.GTS.TRI )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_881 .INIT = 16'h7C4A;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_881  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_88 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_891 .INIT = 16'h43E9;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_891  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_89 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_901 .INIT = 16'hC3A5;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_901  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_90 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_911 .INIT = 16'h9D92;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_911  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[14] ),
    .ADR2(\c1/X[15] ),
    .ADR3(\c1/X[17] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_91 )
  );
  X_BUF key_50_IBUF_125 (
    .I(key[50]),
    .O(key_50_IBUF)
  );
  X_BUF dataout_35_OBUF (
    .I(dataout_35),
    .O(\dataout_35_OBUF.GTS.TRI )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_921 .INIT = 16'h9749;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_921  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[17] ),
    .ADR2(\c1/X[14] ),
    .ADR3(\c1/X[15] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_92 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_931 .INIT = 16'h7AC1;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_931  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[14] ),
    .ADR3(\c1/X[17] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_93 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_941 .INIT = 16'h6693;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_941  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_94 )
  );
  defparam \c1/u2/Mrom_dout_inst_lut4_951 .INIT = 16'h936C;
  X_LUT4 \c1/u2/Mrom_dout_inst_lut4_951  (
    .ADR0(\c1/X[16] ),
    .ADR1(\c1/X[15] ),
    .ADR2(\c1/X[17] ),
    .ADR3(\c1/X[14] ),
    .O(\c1/u2/Mrom_dout_inst_lut4_95 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_961 .INIT = 16'h9E34;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_961  (
    .ADR0(N5937),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_96 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_971 .INIT = 16'h69E2;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_971  (
    .ADR0(N5936),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[4] ),
    .ADR3(\c1/X[2] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_97 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_981 .INIT = 16'h5D92;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_981  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[3] ),
    .ADR2(\c1/X[4] ),
    .ADR3(\c1/X[5] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_98 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_991 .INIT = 16'hA665;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_991  (
    .ADR0(\c1/X[4] ),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[2] ),
    .ADR3(\c1/X[3] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_99 )
  );
  X_BUF dataout_39_OBUF (
    .I(dataout_39),
    .O(\dataout_39_OBUF.GTS.TRI )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1001 .INIT = 16'h8667;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1001  (
    .ADR0(N5939),
    .ADR1(\c1/X[4] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[2] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_100 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1011 .INIT = 16'h3596;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1011  (
    .ADR0(\c1/X[3] ),
    .ADR1(\c1/X[4] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[2] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_101 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1021 .INIT = 16'h3E94;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1021  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_102 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1031 .INIT = 16'h6E49;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1031  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[4] ),
    .ADR3(\c1/X[3] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_103 )
  );
  X_BUF dataout_38_OBUF (
    .I(dataout_38),
    .O(\dataout_38_OBUF.GTS.TRI )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1041 .INIT = 16'h86D3;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1041  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_104 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1051 .INIT = 16'h17A6;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1051  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[4] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[3] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_105 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1061 .INIT = 16'h3497;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1061  (
    .ADR0(\c1/X[3] ),
    .ADR1(\c1/X[4] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[2] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_106 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1071 .INIT = 16'hC993;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1071  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[3] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_107 )
  );
  X_BUF dataout_37_OBUF (
    .I(dataout_37),
    .O(\dataout_37_OBUF.GTS.TRI )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1081 .INIT = 16'h6E31;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1081  (
    .ADR0(N5938),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[2] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_108 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1091 .INIT = 16'hB456;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1091  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[4] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[3] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_109 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1101 .INIT = 16'h297C;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1101  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[3] ),
    .ADR2(\c1/X[5] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_110 )
  );
  defparam \c1/u0/Mrom_dout_inst_lut4_1111 .INIT = 16'h869B;
  X_LUT4 \c1/u0/Mrom_dout_inst_lut4_1111  (
    .ADR0(\c1/X[2] ),
    .ADR1(\c1/X[5] ),
    .ADR2(\c1/X[3] ),
    .ADR3(\c1/X[4] ),
    .O(\c1/u0/Mrom_dout_inst_lut4_111 )
  );
  X_BUF key_47_IBUF_126 (
    .I(key[47]),
    .O(key_47_IBUF)
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1121 .INIT = 16'h2D65;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1121  (
    .ADR0(N5916),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_112 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1131 .INIT = 16'hE21D;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1131  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(N5917),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_113 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1151 .INIT = 16'hC359;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1151  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_115 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_63 .INIT = 16'h8697;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_63  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[11] ),
    .ADR2(N5184),
    .ADR3(N5183),
    .O(\c1/u1/Mrom_dout_N10 )
  );
  X_BUF dataout_30_OBUF (
    .I(dataout_30),
    .O(\dataout_30_OBUF.GTS.TRI )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1171 .INIT = 16'h38D9;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1171  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_117 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1191 .INIT = 16'h27D2;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1191  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_119 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_57 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_57  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_114 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_115 ),
    .O(\c1/u1/Mrom_dout_N1 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_58 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_58  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_116 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_117 ),
    .O(\c1/u1/Mrom_dout_N3 )
  );
  X_BUF dataout_52_OBUF (
    .I(dataout_52),
    .O(\dataout_52_OBUF.GTS.TRI )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1211 .INIT = 16'h919E;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1211  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_121 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1231 .INIT = 16'h6E61;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1231  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_123 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_59 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_59  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_118 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_119 ),
    .O(\c1/u1/Mrom_dout_N4 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_60 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_60  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_120 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_121 ),
    .O(\c1/u1/Mrom_dout_N6 )
  );
  X_BUF dataout_49_OBUF (
    .I(dataout_49),
    .O(\dataout_49_OBUF.GTS.TRI )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_62_SW0 .INIT = 16'h6906;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_62_SW0  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(N5918),
    .ADR3(\c1/X[10] ),
    .O(N5186)
  );
  defparam _n0011_SW0.INIT = 8'hEA;
  X_LUT3 _n0011_SW0 (
    .ADR0(ready_OBUF),
    .ADR1(_n0001),
    .ADR2(state_FFd2),
    .O(N234)
  );
  defparam \_n0012<1>1051_G .INIT = 16'h2882;
  X_LUT4 \_n0012<1>1051_G  (
    .ADR0(rst_IBUF),
    .ADR1(roundsel[1]),
    .ADR2(state_FFd6),
    .ADR3(roundsel[2]),
    .O(N5761)
  );
  defparam \_n0013<39>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<39>8  (
    .ADR0(data1[8]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE785),
    .ADR3(state_FFd5),
    .O(CHOICE787)
  );
  defparam \_n0012<3>33 .INIT = 16'h2878;
  X_LUT4 \_n0012<3>33  (
    .ADR0(_n0025),
    .ADR1(\Maddsub__n0017_Mxor_Result<3>_Xo [0]),
    .ADR2(roundsel[4]),
    .ADR3(state_FFd7),
    .O(CHOICE13)
  );
  defparam \_n0012<3>5 .INIT = 8'hA2;
  X_LUT3 \_n0012<3>5  (
    .ADR0(flag_IBUF),
    .ADR1(rst_IBUF),
    .ADR2(state_FFd7),
    .O(CHOICE2)
  );
  defparam \_n0013<17>6 .INIT = 4'h8;
  X_LUT2 \_n0013<17>6  (
    .ADR0(data1[18]),
    .ADR1(N01),
    .O(CHOICE1047)
  );
  defparam \key2<17>12 .INIT = 16'hCA00;
  X_LUT4 \key2<17>12  (
    .ADR0(\key1[19] ),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_1_10),
    .ADR3(roundsel_23),
    .O(CHOICE521)
  );
  defparam \_n0013<48>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<48>8  (
    .ADR0(data1[17]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE91),
    .ADR3(state_FFd5),
    .O(CHOICE93)
  );
  X_BUF dataout_56_OBUF (
    .I(dataout_56),
    .O(\dataout_56_OBUF.GTS.TRI )
  );
  defparam \_n0013<34>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<34>8  (
    .ADR0(data1[3]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE154),
    .ADR3(state_FFd5),
    .O(CHOICE156)
  );
  defparam \key2<36>74 .INIT = 8'hCA;
  X_LUT3 \key2<36>74  (
    .ADR0(\key1[62] ),
    .ADR1(\key1[5] ),
    .ADR2(roundsel_1_14),
    .O(CHOICE391)
  );
  defparam \_n0013<47>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<47>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[62]),
    .ADR2(state_FFd8),
    .ADR3(datain_48_IBUF),
    .O(CHOICE758)
  );
  defparam \_n0013<30>9 .INIT = 8'hEA;
  X_LUT3 \_n0013<30>9  (
    .ADR0(CHOICE822),
    .ADR1(data1[4]),
    .ADR2(\state_FFd3-In ),
    .O(CHOICE824)
  );
  defparam \_n0013<2>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<2>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[23]),
    .ADR2(state_FFd8),
    .ADR3(datain_3_IBUF),
    .O(CHOICE669)
  );
  defparam \_n0013<42>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<42>8  (
    .ADR0(data1[11]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE19),
    .ADR3(state_FFd5),
    .O(CHOICE21)
  );
  defparam \_n0013<30>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<30>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[49]),
    .ADR2(state_FFd8),
    .ADR3(datain_31_IBUF),
    .O(CHOICE822)
  );
  defparam \_n0012<2>100_SW3 .INIT = 16'hB115;
  X_LUT4 \_n0012<2>100_SW3  (
    .ADR0(state_FFd6),
    .ADR1(state_FFd5),
    .ADR2(roundsel[1]),
    .ADR3(roundsel[2]),
    .O(N5500)
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_61 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_61  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_122 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_123 ),
    .O(\c1/u1/Mrom_dout_N7 )
  );
  defparam \_n0013<1>6 .INIT = 4'h8;
  X_LUT2 \_n0013<1>6  (
    .ADR0(data1[2]),
    .ADR1(N01),
    .O(CHOICE1946)
  );
  X_BUF datain_50_IBUF_127 (
    .I(datain[50]),
    .O(datain_50_IBUF)
  );
  defparam Ker020.INIT = 16'h0001;
  X_LUT4 Ker020 (
    .ADR0(state_FFd8),
    .ADR1(state_FFd7),
    .ADR2(state_FFd5),
    .ADR3(N5428),
    .O(CHOICE195)
  );
  defparam \_n0013<46>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<46>8  (
    .ADR0(data1[15]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE100),
    .ADR3(state_FFd5),
    .O(CHOICE102)
  );
  X_BUF dataout_8_OBUF (
    .I(dataout_8),
    .O(\dataout_8_OBUF.GTS.TRI )
  );
  defparam \_n0013<6>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<6>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[55]),
    .ADR2(state_FFd8),
    .ADR3(datain_7_IBUF),
    .O(CHOICE633)
  );
  defparam \_n0013<49>12 .INIT = 4'h8;
  X_LUT2 \_n0013<49>12  (
    .ADR0(data1[50]),
    .ADR1(N01),
    .O(CHOICE752)
  );
  defparam \_n0013<17>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<17>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[11]),
    .ADR2(state_FFd8),
    .ADR3(datain_18_IBUF),
    .O(CHOICE1046)
  );
  defparam \key2<21>12 .INIT = 16'hCA00;
  X_LUT4 \key2<21>12  (
    .ADR0(\key1[58] ),
    .ADR1(\key1[3] ),
    .ADR2(roundsel_1_10),
    .ADR3(roundsel_2_7),
    .O(CHOICE970)
  );
  defparam \_n0013<32>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<32>8  (
    .ADR0(data1[1]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE145),
    .ADR3(state_FFd5),
    .O(CHOICE147)
  );
  defparam \_n0013<33>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<33>22_SW0  (
    .ADR0(data1[2]),
    .ADR1(_n0025),
    .ADR2(data1[34]),
    .ADR3(N01),
    .O(N5444)
  );
  defparam \_n0013<59>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<59>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[26]),
    .ADR2(state_FFd8),
    .ADR3(datain_60_IBUF),
    .O(CHOICE704)
  );
  X_BUF dataout_10_OBUF (
    .I(dataout_10),
    .O(\dataout_10_OBUF.GTS.TRI )
  );
  defparam \key2<14>74 .INIT = 8'hAC;
  X_LUT3 \key2<14>74  (
    .ADR0(\key1[50] ),
    .ADR1(\key1[42] ),
    .ADR2(roundsel_1_18),
    .O(CHOICE571)
  );
  defparam \_n0013<33>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<33>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[16]),
    .ADR2(state_FFd8),
    .ADR3(datain_34_IBUF),
    .O(CHOICE812)
  );
  defparam \_n0013<62>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<62>8  (
    .ADR0(data1[31]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE28),
    .ADR3(state_FFd5),
    .O(CHOICE30)
  );
  defparam \_n0013<49>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<49>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[12]),
    .ADR2(state_FFd8),
    .ADR3(datain_50_IBUF),
    .O(CHOICE749)
  );
  X_BUF datain_34_IBUF_128 (
    .I(datain[34]),
    .O(datain_34_IBUF)
  );
  defparam Ker030.INIT = 4'h2;
  X_LUT2 Ker030 (
    .ADR0(state_FFd4),
    .ADR1(N5901),
    .O(CHOICE199)
  );
  defparam \_n0013<44>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<44>8  (
    .ADR0(data1[13]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE109),
    .ADR3(state_FFd5),
    .O(CHOICE111)
  );
  defparam \key2<27>97 .INIT = 8'hAC;
  X_LUT3 \key2<27>97  (
    .ADR0(\key1[46] ),
    .ADR1(\key1[38] ),
    .ADR2(roundsel_1_16),
    .O(CHOICE1332)
  );
  X_BUF datain_8_IBUF_129 (
    .I(datain[8]),
    .O(datain_8_IBUF)
  );
  defparam \_n0013<0>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<0>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[7]),
    .ADR2(state_FFd8),
    .ADR3(datain_1_IBUF),
    .O(CHOICE660)
  );
  defparam \_n0013<35>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<35>22_SW0  (
    .ADR0(data1[4]),
    .ADR1(_n0025),
    .ADR2(data1[36]),
    .ADR3(N01),
    .O(N5476)
  );
  defparam \key2<16>61 .INIT = 8'hE4;
  X_LUT3 \key2<16>61  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out62 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out48 ),
    .O(CHOICE510)
  );
  X_BUF dataout_57_OBUF (
    .I(dataout_57),
    .O(\dataout_57_OBUF.GTS.TRI )
  );
  defparam \_n0013<35>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<35>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[32]),
    .ADR2(state_FFd8),
    .ADR3(datain_36_IBUF),
    .O(CHOICE803)
  );
  defparam \_n0013<60>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<60>8  (
    .ADR0(data1[29]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE37),
    .ADR3(state_FFd5),
    .O(CHOICE39)
  );
  defparam \_n0012<2>100 .INIT = 16'h25AD;
  X_LUT4 \_n0012<2>100  (
    .ADR0(roundsel[3]),
    .ADR1(state_FFd7),
    .ADR2(N5499),
    .ADR3(N5500),
    .O(CHOICE230)
  );
  defparam \_n0013<58>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<58>8  (
    .ADR0(data1[27]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE46),
    .ADR3(state_FFd5),
    .O(CHOICE48)
  );
  defparam \_n0013<9>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<9>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[13]),
    .ADR2(state_FFd8),
    .ADR3(datain_10_IBUF),
    .O(CHOICE1927)
  );
  X_BUF datain_30_IBUF_130 (
    .I(datain[30]),
    .O(datain_30_IBUF)
  );
  defparam \_n0013<45>8 .INIT = 8'hA8;
  X_LUT3 \_n0013<45>8  (
    .ADR0(data1[46]),
    .ADR1(state_FFd7),
    .ADR2(N01),
    .O(CHOICE626)
  );
  defparam \_n0013<61>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<61>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[42]),
    .ADR2(state_FFd8),
    .ADR3(datain_62_IBUF),
    .O(CHOICE695)
  );
  defparam \_n0013<51>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<51>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[28]),
    .ADR2(state_FFd8),
    .ADR3(datain_52_IBUF),
    .O(CHOICE740)
  );
  X_BUF datain_49_IBUF_131 (
    .I(datain[49]),
    .O(datain_49_IBUF)
  );
  X_BUF dataout_7_OBUF (
    .I(dataout_7),
    .O(\dataout_7_OBUF.GTS.TRI )
  );
  X_BUF dataout_1_OBUF (
    .I(dataout_1),
    .O(\dataout_1_OBUF.GTS.TRI )
  );
  defparam \_n0013<45>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<45>5  (
    .ADR0(state_FFd8),
    .ADR1(datain_46_IBUF),
    .ADR2(data1[14]),
    .ADR3(_n0025),
    .O(CHOICE624)
  );
  defparam \_n0013<40>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<40>8  (
    .ADR0(data1[9]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE118),
    .ADR3(state_FFd5),
    .O(CHOICE120)
  );
  X_BUF dataout_61_OBUF (
    .I(dataout_61),
    .O(\dataout_61_OBUF.GTS.TRI )
  );
  defparam \_n0013<37>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<37>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[48]),
    .ADR2(state_FFd8),
    .ADR3(datain_38_IBUF),
    .O(CHOICE794)
  );
  defparam \key2<24>74 .INIT = 8'hE4;
  X_LUT3 \key2<24>74  (
    .ADR0(roundsel[1]),
    .ADR1(\key1[43] ),
    .ADR2(\key1[51] ),
    .O(CHOICE423)
  );
  defparam roundsel_2_8_132.INIT = 1'b1;
  X_SFF roundsel_2_8_132 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_8),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  X_BUF dataout_63_OBUF (
    .I(dataout_63),
    .O(\dataout_63_OBUF.GTS.TRI )
  );
  defparam \_n0013<54>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<54>8  (
    .ADR0(data1[23]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE55),
    .ADR3(state_FFd5),
    .O(CHOICE57)
  );
  defparam \_n0013<53>12 .INIT = 4'h8;
  X_LUT2 \_n0013<53>12  (
    .ADR0(data1[54]),
    .ADR1(N01),
    .O(CHOICE734)
  );
  defparam \_n0013<49>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<49>8  (
    .ADR0(data1[18]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE749),
    .ADR3(state_FFd5),
    .O(CHOICE751)
  );
  defparam \_n0013<1>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<1>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[15]),
    .ADR2(state_FFd8),
    .ADR3(datain_2_IBUF),
    .O(CHOICE1945)
  );
  defparam \_n0013<63>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<63>22_SW0  (
    .ADR0(data1[32]),
    .ADR1(_n0025),
    .ADR2(data1[64]),
    .ADR3(N01),
    .O(N5460)
  );
  defparam \_n0013<10>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<10>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[21]),
    .ADR2(state_FFd8),
    .ADR3(datain_11_IBUF),
    .O(CHOICE651)
  );
  defparam \_n0013<38>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<38>8  (
    .ADR0(data1[7]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE127),
    .ADR3(state_FFd5),
    .O(CHOICE129)
  );
  defparam \_n0013<53>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<53>8  (
    .ADR0(data1[22]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE731),
    .ADR3(state_FFd5),
    .O(CHOICE733)
  );
  defparam \_n0013<53>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<53>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[44]),
    .ADR2(state_FFd8),
    .ADR3(datain_54_IBUF),
    .O(CHOICE731)
  );
  X_BUF dataout_62_OBUF (
    .I(dataout_62),
    .O(\dataout_62_OBUF.GTS.TRI )
  );
  defparam \_n0013<63>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<63>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[58]),
    .ADR2(state_FFd8),
    .ADR3(datain_64_IBUF),
    .O(CHOICE686)
  );
  defparam \_n0013<39>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<39>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[64]),
    .ADR2(state_FFd8),
    .ADR3(datain_40_IBUF),
    .O(CHOICE785)
  );
  defparam \key2<1>61 .INIT = 8'hE4;
  X_LUT3 \key2<1>61  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out75 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out29 ),
    .O(CHOICE1093)
  );
  defparam \_n0013<9>6 .INIT = 4'h8;
  X_LUT2 \_n0013<9>6  (
    .ADR0(data1[10]),
    .ADR1(N01),
    .O(CHOICE1928)
  );
  X_BUF datain_9_IBUF_133 (
    .I(datain[9]),
    .O(datain_9_IBUF)
  );
  defparam \_n0013<56>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<56>8  (
    .ADR0(data1[25]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE64),
    .ADR3(state_FFd5),
    .O(CHOICE66)
  );
  X_BUF datain_51_IBUF_134 (
    .I(datain[51]),
    .O(datain_51_IBUF)
  );
  defparam \_n0013<36>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<36>8  (
    .ADR0(data1[5]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE136),
    .ADR3(state_FFd5),
    .O(CHOICE138)
  );
  defparam \_n0013<18>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<18>5  (
    .ADR0(state_FFd8),
    .ADR1(datain_19_IBUF),
    .ADR2(data1[19]),
    .ADR3(\state_FFd3-In ),
    .O(CHOICE616)
  );
  defparam \_n0013<41>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<41>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[14]),
    .ADR2(state_FFd8),
    .ADR3(datain_42_IBUF),
    .O(CHOICE776)
  );
  defparam \_n0013<55>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<55>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[60]),
    .ADR2(state_FFd8),
    .ADR3(datain_56_IBUF),
    .O(CHOICE722)
  );
  defparam \_n0013<4>9 .INIT = 8'hEA;
  X_LUT3 \_n0013<4>9  (
    .ADR0(CHOICE678),
    .ADR1(data1[9]),
    .ADR2(\state_FFd3-In ),
    .O(CHOICE680)
  );
  defparam \key2<30>74 .INIT = 8'hAC;
  X_LUT3 \key2<30>74  (
    .ADR0(\key1[14] ),
    .ADR1(\key1[6] ),
    .ADR2(roundsel_1_14),
    .O(CHOICE455)
  );
  X_BUF datain_48_IBUF_135 (
    .I(datain[48]),
    .O(datain_48_IBUF)
  );
  defparam \_n0013<4>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<4>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[39]),
    .ADR2(state_FFd8),
    .ADR3(datain_5_IBUF),
    .O(CHOICE678)
  );
  defparam \_n0013<52>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<52>8  (
    .ADR0(data1[21]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE73),
    .ADR3(state_FFd5),
    .O(CHOICE75)
  );
  X_BUF dataout_64_OBUF (
    .I(dataout_64),
    .O(\dataout_64_OBUF.GTS.TRI )
  );
  defparam \key2<16>12 .INIT = 16'hA280;
  X_LUT4 \key2<16>12  (
    .ADR0(roundsel_2_6),
    .ADR1(roundsel_3_11),
    .ADR2(N5905),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out52 ),
    .O(CHOICE497)
  );
  defparam \_n0013<50>8 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<50>8  (
    .ADR0(data1[19]),
    .ADR1(state_FFd6),
    .ADR2(CHOICE82),
    .ADR3(state_FFd5),
    .O(CHOICE84)
  );
  defparam \_n0013<8>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<8>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[5]),
    .ADR2(state_FFd8),
    .ADR3(datain_9_IBUF),
    .O(CHOICE642)
  );
  X_BUF dataout_11_OBUF (
    .I(dataout_11),
    .O(\dataout_11_OBUF.GTS.TRI )
  );
  defparam \_n0013<43>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<43>22_SW0  (
    .ADR0(data1[12]),
    .ADR1(_n0025),
    .ADR2(data1[44]),
    .ADR3(N01),
    .O(N5442)
  );
  defparam \_n0013<4>1 .INIT = 4'h8;
  X_LUT2 \_n0013<4>1  (
    .ADR0(data1[5]),
    .ADR1(N5900),
    .O(CHOICE675)
  );
  defparam \_n0013<43>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<43>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[30]),
    .ADR2(state_FFd8),
    .ADR3(datain_44_IBUF),
    .O(CHOICE767)
  );
  defparam \key2<15>25_SW0 .INIT = 16'hFF53;
  X_LUT4 \key2<15>25_SW0  (
    .ADR0(\key1[43] ),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_22),
    .O(N5129)
  );
  X_BUF datain_26_IBUF_136 (
    .I(datain[26]),
    .O(datain_26_IBUF)
  );
  X_BUF datain_11_IBUF_137 (
    .I(datain[11]),
    .O(datain_11_IBUF)
  );
  X_BUF key_2_IBUF_138 (
    .I(key[2]),
    .O(key_2_IBUF)
  );
  defparam \_n0013<7>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<7>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[63]),
    .ADR2(state_FFd8),
    .ADR3(datain_8_IBUF),
    .O(CHOICE1918)
  );
  X_BUF key_55_IBUF_139 (
    .I(key[55]),
    .O(key_55_IBUF)
  );
  X_BUF key_12_IBUF_140 (
    .I(key[12]),
    .O(key_12_IBUF)
  );
  defparam \key2<3>74 .INIT = 8'hAC;
  X_LUT3 \key2<3>74  (
    .ADR0(\key1[11] ),
    .ADR1(\key1[3] ),
    .ADR2(roundsel_1_18),
    .O(CHOICE1577)
  );
  defparam \_n0013<26>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<26>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[17]),
    .ADR2(state_FFd8),
    .ADR3(datain_27_IBUF),
    .O(CHOICE840)
  );
  X_BUF key_46_IBUF_141 (
    .I(key[46]),
    .O(key_46_IBUF)
  );
  X_BUF dataout_12_OBUF (
    .I(dataout_12),
    .O(\dataout_12_OBUF.GTS.TRI )
  );
  defparam \_n0013<29>6 .INIT = 4'h8;
  X_LUT2 \_n0013<29>6  (
    .ADR0(data1[30]),
    .ADR1(N01),
    .O(CHOICE1955)
  );
  X_BUF key_37_IBUF_142 (
    .I(key[37]),
    .O(key_37_IBUF)
  );
  X_BUF key_60_IBUF_143 (
    .I(key[60]),
    .O(key_60_IBUF)
  );
  X_BUF key_19_IBUF_144 (
    .I(key[19]),
    .O(key_19_IBUF)
  );
  defparam \key2<45>12 .INIT = 16'hCA00;
  X_LUT4 \key2<45>12  (
    .ADR0(\key1[54] ),
    .ADR1(\key1[62] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_2_1),
    .O(CHOICE1855)
  );
  X_BUF datain_28_IBUF_145 (
    .I(datain[28]),
    .O(datain_28_IBUF)
  );
  defparam \_n0013<15>6 .INIT = 4'h8;
  X_LUT2 \_n0013<15>6  (
    .ADR0(data1[16]),
    .ADR1(N01),
    .O(CHOICE2009)
  );
  defparam \_n0013<15>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<15>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[61]),
    .ADR2(state_FFd8),
    .ADR3(datain_16_IBUF),
    .O(CHOICE2008)
  );
  X_BUF key_4_IBUF_146 (
    .I(key[4]),
    .O(key_4_IBUF)
  );
  X_BUF key_6_IBUF_147 (
    .I(key[6]),
    .O(key_6_IBUF)
  );
  X_BUF datain_14_IBUF_148 (
    .I(datain[14]),
    .O(datain_14_IBUF)
  );
  X_BUF key_8_IBUF_149 (
    .I(key[8]),
    .O(key_8_IBUF)
  );
  X_BUF key_32_IBUF_150 (
    .I(key[32]),
    .O(key_32_IBUF)
  );
  X_BUF datain_13_IBUF_151 (
    .I(datain[13]),
    .O(datain_13_IBUF)
  );
  X_BUF key_56_IBUF_152 (
    .I(key[56]),
    .O(key_56_IBUF)
  );
  X_BUF datain_20_IBUF_153 (
    .I(datain[20]),
    .O(datain_20_IBUF)
  );
  X_BUF key_34_IBUF_154 (
    .I(key[34]),
    .O(key_34_IBUF)
  );
  defparam \key2<19>15 .INIT = 16'h0E04;
  X_LUT4 \key2<19>15  (
    .ADR0(roundsel[2]),
    .ADR1(N5903),
    .ADR2(roundsel[3]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out38 ),
    .O(CHOICE851)
  );
  X_BUF key_51_IBUF_155 (
    .I(key[51]),
    .O(key_51_IBUF)
  );
  defparam \_n0013<22>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<22>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[51]),
    .ADR2(state_FFd8),
    .ADR3(datain_23_IBUF),
    .O(CHOICE1020)
  );
  X_BUF dataout_19_OBUF (
    .I(dataout_19),
    .O(\dataout_19_OBUF.GTS.TRI )
  );
  defparam \_n0013<29>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<29>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[41]),
    .ADR2(state_FFd8),
    .ADR3(datain_30_IBUF),
    .O(CHOICE1954)
  );
  X_BUF key_11_IBUF_156 (
    .I(key[11]),
    .O(key_11_IBUF)
  );
  defparam \_n0013<31>6 .INIT = 4'h8;
  X_LUT2 \_n0013<31>6  (
    .ADR0(data1[32]),
    .ADR1(Ker039),
    .O(CHOICE1964)
  );
  defparam \key2<45>25_SW0 .INIT = 16'hFF53;
  X_LUT4 \key2<45>25_SW0  (
    .ADR0(\key1[38] ),
    .ADR1(\key1[22] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_22),
    .O(N5137)
  );
  defparam \_n0013<19>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<19>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[27]),
    .ADR2(state_FFd8),
    .ADR3(datain_20_IBUF),
    .O(CHOICE1999)
  );
  X_BUF datain_40_IBUF_157 (
    .I(datain[40]),
    .O(datain_40_IBUF)
  );
  X_BUF key_13_IBUF_158 (
    .I(key[13]),
    .O(key_13_IBUF)
  );
  X_BUF key_15_IBUF_159 (
    .I(key[15]),
    .O(key_15_IBUF)
  );
  X_BUF key_18_IBUF_160 (
    .I(key[18]),
    .O(key_18_IBUF)
  );
  X_BUF key_54_IBUF_161 (
    .I(key[54]),
    .O(key_54_IBUF)
  );
  X_BUF key_20_IBUF_162 (
    .I(key[20]),
    .O(key_20_IBUF)
  );
  defparam \_n0013<31>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<31>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[57]),
    .ADR2(state_FFd8),
    .ADR3(datain_32_IBUF),
    .O(CHOICE1963)
  );
  defparam \key2<46>25_SW0 .INIT = 16'hF5F3;
  X_LUT4 \key2<46>25_SW0  (
    .ADR0(\key1[32] ),
    .ADR1(\key1[16] ),
    .ADR2(roundsel_32),
    .ADR3(roundsel_12),
    .O(N5139)
  );
  X_BUF datain_64_IBUF_163 (
    .I(datain[64]),
    .O(datain_64_IBUF)
  );
  X_BUF datain_46_IBUF_164 (
    .I(datain[46]),
    .O(datain_46_IBUF)
  );
  X_BUF dataout_22_OBUF (
    .I(dataout_22),
    .O(\dataout_22_OBUF.GTS.TRI )
  );
  X_BUF rst_IBUF_165 (
    .I(rst),
    .O(rst_IBUF)
  );
  defparam \_n0013<24>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<24>22_SW0  (
    .ADR0(data1[28]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[25]),
    .ADR3(N01),
    .O(N5480)
  );
  X_BUF key_3_IBUF_166 (
    .I(key[3]),
    .O(key_3_IBUF)
  );
  X_BUF datain_16_IBUF_167 (
    .I(datain[16]),
    .O(datain_16_IBUF)
  );
  X_BUF datain_44_IBUF_168 (
    .I(datain[44]),
    .O(datain_44_IBUF)
  );
  X_BUF key_26_IBUF_169 (
    .I(key[26]),
    .O(key_26_IBUF)
  );
  X_BUF key_38_IBUF_170 (
    .I(key[38]),
    .O(key_38_IBUF)
  );
  X_BUF dataout_59_OBUF (
    .I(dataout_59),
    .O(\dataout_59_OBUF.GTS.TRI )
  );
  defparam \_n0013<23>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<23>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[59]),
    .ADR2(state_FFd8),
    .ADR3(datain_24_IBUF),
    .O(CHOICE1276)
  );
  X_BUF key_44_IBUF_171 (
    .I(key[44]),
    .O(key_44_IBUF)
  );
  defparam \_n0013<21>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<21>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[43]),
    .ADR2(state_FFd8),
    .ADR3(datain_22_IBUF),
    .O(CHOICE1990)
  );
  defparam \_n0013<24>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<24>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[1]),
    .ADR2(state_FFd8),
    .ADR3(datain_25_IBUF),
    .O(CHOICE1002)
  );
  X_BUF key_16_IBUF_172 (
    .I(key[16]),
    .O(key_16_IBUF)
  );
  defparam \_n0013<5>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<5>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[47]),
    .ADR2(state_FFd8),
    .ADR3(datain_6_IBUF),
    .O(CHOICE1267)
  );
  X_BUF datain_24_IBUF_173 (
    .I(datain[24]),
    .O(datain_24_IBUF)
  );
  defparam \_n0013<5>6 .INIT = 4'h8;
  X_LUT2 \_n0013<5>6  (
    .ADR0(data1[6]),
    .ADR1(N01),
    .O(CHOICE1268)
  );
  defparam \_n0013<12>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<12>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[37]),
    .ADR2(state_FFd8),
    .ADR3(datain_13_IBUF),
    .O(CHOICE1029)
  );
  X_BUF datain_52_IBUF_174 (
    .I(datain[52]),
    .O(datain_52_IBUF)
  );
  X_BUF dataout_20_OBUF (
    .I(dataout_20),
    .O(\dataout_20_OBUF.GTS.TRI )
  );
  X_BUF datain_36_IBUF_175 (
    .I(datain[36]),
    .O(datain_36_IBUF)
  );
  X_BUF key_21_IBUF_176 (
    .I(key[21]),
    .O(key_21_IBUF)
  );
  defparam \_n0013<23>6 .INIT = 4'h8;
  X_LUT2 \_n0013<23>6  (
    .ADR0(data1[24]),
    .ADR1(N01),
    .O(CHOICE1277)
  );
  X_BUF key_30_IBUF_177 (
    .I(key[30]),
    .O(key_30_IBUF)
  );
  X_BUF key_58_IBUF_178 (
    .I(key[58]),
    .O(key_58_IBUF)
  );
  defparam \key2<27>12 .INIT = 16'hAC00;
  X_LUT4 \key2<27>12  (
    .ADR0(\key1[30] ),
    .ADR1(\key1[22] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_3_1),
    .O(CHOICE1310)
  );
  X_BUF dataout_16_OBUF (
    .I(dataout_16),
    .O(\dataout_16_OBUF.GTS.TRI )
  );
  X_BUF key_22_IBUF_179 (
    .I(key[22]),
    .O(key_22_IBUF)
  );
  X_BUF datain_42_IBUF_180 (
    .I(datain[42]),
    .O(datain_42_IBUF)
  );
  X_BUF datain_15_IBUF_181 (
    .I(datain[15]),
    .O(datain_15_IBUF)
  );
  X_BUF datain_17_IBUF_182 (
    .I(datain[17]),
    .O(datain_17_IBUF)
  );
  X_BUF datain_18_IBUF_183 (
    .I(datain[18]),
    .O(datain_18_IBUF)
  );
  defparam \_n0013<25>6 .INIT = 4'h8;
  X_LUT2 \_n0013<25>6  (
    .ADR0(data1[26]),
    .ADR1(N01),
    .O(CHOICE1982)
  );
  defparam \_n0013<25>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<25>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[9]),
    .ADR2(state_FFd8),
    .ADR3(datain_26_IBUF),
    .O(CHOICE1981)
  );
  X_BUF dataout_23_OBUF (
    .I(dataout_23),
    .O(\dataout_23_OBUF.GTS.TRI )
  );
  X_BUF key_14_IBUF_184 (
    .I(key[14]),
    .O(key_14_IBUF)
  );
  X_BUF datain_55_IBUF_185 (
    .I(datain[55]),
    .O(datain_55_IBUF)
  );
  X_BUF dataout_14_OBUF (
    .I(dataout_14),
    .O(\dataout_14_OBUF.GTS.TRI )
  );
  X_BUF key_10_IBUF_186 (
    .I(key[10]),
    .O(key_10_IBUF)
  );
  X_BUF datain_54_IBUF_187 (
    .I(datain[54]),
    .O(datain_54_IBUF)
  );
  defparam \_n0013<16>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<16>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[3]),
    .ADR2(state_FFd8),
    .ADR3(datain_17_IBUF),
    .O(CHOICE873)
  );
  X_BUF datain_62_IBUF_188 (
    .I(datain[62]),
    .O(datain_62_IBUF)
  );
  defparam \_n0013<20>6 .INIT = 16'hF888;
  X_LUT4 \_n0013<20>6  (
    .ADR0(state_FFd7),
    .ADR1(data1[35]),
    .ADR2(state_FFd8),
    .ADR3(datain_21_IBUF),
    .O(CHOICE1011)
  );
  X_BUF dataout_15_OBUF (
    .I(dataout_15),
    .O(\dataout_15_OBUF.GTS.TRI )
  );
  X_BUF key_24_IBUF_189 (
    .I(key[24]),
    .O(key_24_IBUF)
  );
  defparam \key2<1>12 .INIT = 16'hA280;
  X_LUT4 \key2<1>12  (
    .ADR0(roundsel[2]),
    .ADR1(roundsel[3]),
    .ADR2(N5904),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out47 ),
    .O(CHOICE1080)
  );
  defparam \key2<23>74 .INIT = 8'hAC;
  X_LUT3 \key2<23>74  (
    .ADR0(\key1[45] ),
    .ADR1(\key1[37] ),
    .ADR2(roundsel_1_9),
    .O(CHOICE900)
  );
  X_BUF key_36_IBUF_190 (
    .I(key[36]),
    .O(key_36_IBUF)
  );
  defparam \key2<32>61 .INIT = 8'hE4;
  X_LUT3 \key2<32>61  (
    .ADR0(roundsel_2_4),
    .ADR1(N5906),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out87 ),
    .O(CHOICE1676)
  );
  X_BUF key_23_IBUF_191 (
    .I(key[23]),
    .O(key_23_IBUF)
  );
  defparam \key2<29>74 .INIT = 8'hAC;
  X_LUT3 \key2<29>74  (
    .ADR0(\key1[7] ),
    .ADR1(\key1[64] ),
    .ADR2(roundsel_1_16),
    .O(CHOICE1545)
  );
  defparam \_n0013<27>6 .INIT = 4'h8;
  X_LUT2 \_n0013<27>6  (
    .ADR0(data1[28]),
    .ADR1(N01),
    .O(CHOICE1973)
  );
  X_BUF dataout_54_OBUF (
    .I(dataout_54),
    .O(\dataout_54_OBUF.GTS.TRI )
  );
  defparam \_n0013<27>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<27>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[25]),
    .ADR2(state_FFd8),
    .ADR3(datain_28_IBUF),
    .O(CHOICE1972)
  );
  defparam \key2<21>25_SW0 .INIT = 16'hFF53;
  X_LUT4 \key2<21>25_SW0  (
    .ADR0(\key1[42] ),
    .ADR1(\key1[26] ),
    .ADR2(roundsel_1_10),
    .ADR3(roundsel_22),
    .O(N5131)
  );
  X_BUF key_53_IBUF_192 (
    .I(key[53]),
    .O(key_53_IBUF)
  );
  X_BUF key_27_IBUF_193 (
    .I(key[27]),
    .O(key_27_IBUF)
  );
  X_BUF datain_53_IBUF_194 (
    .I(datain[53]),
    .O(datain_53_IBUF)
  );
  X_BUF key_29_IBUF_195 (
    .I(key[29]),
    .O(key_29_IBUF)
  );
  X_BUF dataout_18_OBUF (
    .I(dataout_18),
    .O(\dataout_18_OBUF.GTS.TRI )
  );
  X_BUF dataout_13_OBUF (
    .I(dataout_13),
    .O(\dataout_13_OBUF.GTS.TRI )
  );
  X_BUF key_40_IBUF_196 (
    .I(key[40]),
    .O(key_40_IBUF)
  );
  X_BUF datain_32_IBUF_197 (
    .I(datain[32]),
    .O(datain_32_IBUF)
  );
  X_BUF key_31_IBUF_198 (
    .I(key[31]),
    .O(key_31_IBUF)
  );
  defparam roundsel_1_1_199.INIT = 1'b0;
  X_FF roundsel_1_1_199 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_11),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3_1_200.INIT = 1'b1;
  X_SFF roundsel_3_1_200 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_1),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_1_201.INIT = 1'b1;
  X_SFF roundsel_2_1_201 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_1),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_1_202.INIT = 1'b1;
  X_SFF roundsel_4_1_202 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_1),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_2_203.INIT = 1'b0;
  X_FF roundsel_1_2_203 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_1),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3_2_204.INIT = 1'b1;
  X_SFF roundsel_3_2_204 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_32),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_2.INIT = 1'b1;
  X_SFF roundsel_2_2 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_22),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_3_205.INIT = 1'b0;
  X_FF roundsel_1_3_205 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_12),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_4_206.INIT = 1'b0;
  X_FF roundsel_1_4_206 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_11),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_5_207.INIT = 1'b0;
  X_FF roundsel_1_5_207 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_3),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_6_208.INIT = 1'b0;
  X_FF roundsel_1_6_208 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_6),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_2_3.INIT = 1'b1;
  X_SFF roundsel_2_3 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_23),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_3_209.INIT = 1'b1;
  X_SFF roundsel_3_3_209 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_33),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_3_210.INIT = 1'b1;
  X_SFF roundsel_4_3_210 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_43),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_4_211.INIT = 1'b1;
  X_SFF roundsel_2_4_211 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_4),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_7_212.INIT = 1'b0;
  X_FF roundsel_1_7_212 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_2),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_8_213.INIT = 1'b0;
  X_FF roundsel_1_8_213 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_4),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_9_214.INIT = 1'b0;
  X_FF roundsel_1_9_214 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_5),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_10_215.INIT = 1'b0;
  X_FF roundsel_1_10_215 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_10),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3_5_216.INIT = 1'b1;
  X_SFF roundsel_3_5_216 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_3),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_4.INIT = 1'b1;
  X_SFF roundsel_4_4 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_3),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_5_217.INIT = 1'b1;
  X_SFF roundsel_2_5_217 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_24),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_5_218.INIT = 1'b1;
  X_SFF roundsel_4_5_218 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_5),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_6_219.INIT = 1'b1;
  X_SFF roundsel_3_6_219 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_6),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_6_220.INIT = 1'b1;
  X_SFF roundsel_2_6_220 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_6),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_7_221.INIT = 1'b1;
  X_SFF roundsel_2_7_221 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_7),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_7_222.INIT = 1'b1;
  X_SFF roundsel_3_7_222 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_7),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_8_223.INIT = 1'b1;
  X_SFF roundsel_3_8_223 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_8),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_11_224.INIT = 1'b0;
  X_FF roundsel_1_11_224 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_7),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_12.INIT = 1'b0;
  X_FF roundsel_1_12 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_8),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_13.INIT = 1'b0;
  X_FF roundsel_1_13 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_9),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_3_9.INIT = 1'b1;
  X_SFF roundsel_3_9 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_5),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_9.INIT = 1'b1;
  X_SFF roundsel_2_9 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_5),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_10_225.INIT = 1'b1;
  X_SFF roundsel_2_10_225 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_10),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_14_226.INIT = 1'b0;
  X_FF roundsel_1_14_226 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_14),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_4_6_227.INIT = 1'b1;
  X_SFF roundsel_4_6_227 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_6),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_7_228.INIT = 1'b1;
  X_SFF roundsel_4_7_228 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_7),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_8_229.INIT = 1'b1;
  X_SFF roundsel_4_8_229 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_8),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_4_9_230.INIT = 1'b1;
  X_SFF roundsel_4_9_230 (
    .I(N5008),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_4_9),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_10_231.INIT = 1'b1;
  X_SFF roundsel_3_10_231 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_10),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_11_232.INIT = 1'b1;
  X_SFF roundsel_3_11_232 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_11),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_12_233.INIT = 1'b1;
  X_SFF roundsel_3_12_233 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_12),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_13_234.INIT = 1'b1;
  X_SFF roundsel_3_13_234 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_13),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_14_235.INIT = 1'b1;
  X_SFF roundsel_3_14_235 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_14),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_3_15_236.INIT = 1'b1;
  X_SFF roundsel_3_15_236 (
    .I(N5010),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_3_15),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_15_237.INIT = 1'b0;
  X_FF roundsel_1_15_237 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_15),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_16_238.INIT = 1'b0;
  X_FF roundsel_1_16_238 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_16),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_17_239.INIT = 1'b0;
  X_FF roundsel_1_17_239 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_17),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_18_240.INIT = 1'b0;
  X_FF roundsel_1_18_240 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_18),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_19_241.INIT = 1'b0;
  X_FF roundsel_1_19_241 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_19),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_2_11_242.INIT = 1'b1;
  X_SFF roundsel_2_11_242 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_11),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_12_243.INIT = 1'b1;
  X_SFF roundsel_2_12_243 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_12),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_2_13_244.INIT = 1'b1;
  X_SFF roundsel_2_13_244 (
    .I(N5009),
    .SSET(CHOICE2),
    .CLK(clk_BUFGP),
    .O(roundsel_2_13),
    .CE(VCC),
    .SET(GSR),
    .RST(GND),
    .SRST(GND)
  );
  defparam roundsel_1_20_245.INIT = 1'b0;
  X_FF roundsel_1_20_245 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_20),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_21_246.INIT = 1'b0;
  X_FF roundsel_1_21_246 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_21),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam roundsel_1_22_247.INIT = 1'b0;
  X_FF roundsel_1_22_247 (
    .I(_n0012[0]),
    .CLK(clk_BUFGP),
    .O(roundsel_1_22),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  X_MUX2 \key2<22>110_SW01  (
    .IA(N5620),
    .IB(N5621),
    .SEL(roundsel_2_12),
    .O(N5067)
  );
  X_MUX2 \key2<4>110_SW01  (
    .IA(N5622),
    .IB(N5623),
    .SEL(roundsel_2_8),
    .O(N5089)
  );
  X_MUX2 \key2<3>1181  (
    .IA(N5624),
    .IB(N5625),
    .SEL(roundsel_3_3),
    .O(CHOICE1585)
  );
  X_MUX2 \key2<32>271  (
    .IA(N5626),
    .IB(N5627),
    .SEL(roundsel_1_9),
    .O(CHOICE1669)
  );
  X_MUX2 \key2<47>110_SW01  (
    .IA(N5628),
    .IB(N5629),
    .SEL(roundsel_2_11),
    .O(N5083)
  );
  X_MUX2 \key2<28>1191  (
    .IA(N5630),
    .IB(N5631),
    .SEL(roundsel_4_8),
    .O(CHOICE1849)
  );
  X_MUX2 \_n0012<0>  (
    .IA(N5632),
    .IB(N5633),
    .SEL(_n0025),
    .O(_n0012[0])
  );
  defparam \_n0012<0>_F .INIT = 16'hB8AA;
  X_LUT4 \_n0012<0>_F  (
    .ADR0(flag_IBUF),
    .ADR1(state_FFd7),
    .ADR2(roundsel[1]),
    .ADR3(rst_IBUF),
    .O(N5632)
  );
  X_MUX2 \key2<25>961  (
    .IA(N5634),
    .IB(N5635),
    .SEL(roundsel_2_13),
    .O(CHOICE1150)
  );
  X_MUX2 \key2<37>961  (
    .IA(N5636),
    .IB(N5637),
    .SEL(roundsel[2]),
    .O(CHOICE1178)
  );
  X_MUX2 \key2<38>961  (
    .IA(N5638),
    .IB(N5639),
    .SEL(roundsel_2_8),
    .O(CHOICE1817)
  );
  X_MUX2 \key2<3>133_SW01  (
    .IA(N5640),
    .IB(N5641),
    .SEL(roundsel_3_15),
    .O(N5085)
  );
  X_MUX2 \key2<25>12_SW0  (
    .IA(N5642),
    .IB(N5643),
    .SEL(roundsel_3_5),
    .O(N5173)
  );
  X_MUX2 \key2<21>1191  (
    .IA(N5644),
    .IB(N5645),
    .SEL(roundsel_4_5),
    .O(CHOICE996)
  );
  X_MUX2 \key2<33>961  (
    .IA(N5646),
    .IB(N5647),
    .SEL(roundsel_2_4),
    .O(CHOICE1493)
  );
  X_MUX2 \roundsel<2>_mmx_out271  (
    .IA(N5648),
    .IB(N5649),
    .SEL(roundsel_23),
    .O(\MUX_BLOCK_roundsel<2>_mmx_out27 )
  );
  X_MUX2 \key2<22>961  (
    .IA(N5650),
    .IB(N5651),
    .SEL(roundsel_2_12),
    .O(CHOICE936)
  );
  X_MUX2 \key2<32>12  (
    .IA(N5652),
    .IB(N5653),
    .SEL(roundsel_3_2),
    .O(CHOICE1663)
  );
  X_MUX2 \roundsel<2>_mmx_out71  (
    .IA(N5654),
    .IB(N5655),
    .SEL(roundsel_2_7),
    .O(\MUX_BLOCK_roundsel<2>_mmx_out7 )
  );
  X_MUX2 \key2<29>133_SW01  (
    .IA(N5656),
    .IB(N5657),
    .SEL(roundsel_2_5),
    .O(N5071)
  );
  X_MUX2 \key2<41>961  (
    .IA(N5658),
    .IB(N5659),
    .SEL(roundsel_2_5),
    .O(CHOICE1465)
  );
  X_MUX2 \key2<19>761  (
    .IA(N5660),
    .IB(N5661),
    .SEL(roundsel[2]),
    .O(CHOICE867)
  );
  X_MUX2 \roundsel<2>_mmx_out111  (
    .IA(N5662),
    .IB(N5663),
    .SEL(roundsel_2_4),
    .O(\MUX_BLOCK_roundsel<2>_mmx_out11 )
  );
  X_MUX2 \key2<39>761  (
    .IA(N5664),
    .IB(N5665),
    .SEL(roundsel_2_12),
    .O(CHOICE1609)
  );
  X_MUX2 \key2<31>761  (
    .IA(N5666),
    .IB(N5667),
    .SEL(roundsel_24),
    .O(CHOICE1122)
  );
  X_MUX2 \key2<4>961  (
    .IA(N5668),
    .IB(N5669),
    .SEL(roundsel_2_5),
    .O(CHOICE1761)
  );
  X_MUX2 \key2<47>961  (
    .IA(N5670),
    .IB(N5671),
    .SEL(roundsel_2_8),
    .O(CHOICE1377)
  );
  X_MUX2 \key2<44>110_SW01  (
    .IA(N5672),
    .IB(N5673),
    .SEL(roundsel_2_11),
    .O(N5081)
  );
  X_MUX2 \key2<34>110_SW01  (
    .IA(N5674),
    .IB(N5675),
    .SEL(roundsel_22),
    .O(N5075)
  );
  X_MUX2 \key2<43>961  (
    .IA(N5676),
    .IB(N5677),
    .SEL(roundsel[2]),
    .O(CHOICE1206)
  );
  X_MUX2 \c1/Mxor_X_Result<7>11  (
    .IA(N5678),
    .IB(N5679),
    .SEL(roundsel[4]),
    .O(\c1/X[8] )
  );
  X_MUX2 \key2<35>761  (
    .IA(N5680),
    .IB(N5681),
    .SEL(roundsel_2_4),
    .O(CHOICE1304)
  );
  X_MUX2 \key2<45>471  (
    .IA(N5682),
    .IB(N5683),
    .SEL(roundsel_1_22),
    .O(CHOICE1865)
  );
  X_MUX2 \key2<6>110_SW01  (
    .IA(N5684),
    .IB(N5685),
    .SEL(roundsel[2]),
    .O(N5153)
  );
  X_MUX2 \key2<34>961  (
    .IA(N5686),
    .IB(N5687),
    .SEL(roundsel_23),
    .O(CHOICE1234)
  );
  X_MUX2 \key2<6>961  (
    .IA(N5688),
    .IB(N5689),
    .SEL(roundsel[2]),
    .O(CHOICE339)
  );
  X_MUX2 \key2<35>90_SW01  (
    .IA(N5690),
    .IB(N5691),
    .SEL(roundsel_22),
    .O(N5105)
  );
  X_MUX2 \key2<30>1181  (
    .IA(N5692),
    .IB(N5693),
    .SEL(roundsel[2]),
    .O(CHOICE463)
  );
  X_MUX2 \key2<17>471  (
    .IA(N5694),
    .IB(N5695),
    .SEL(roundsel_1_6),
    .O(CHOICE531)
  );
  X_MUX2 \key2<18>961  (
    .IA(N5696),
    .IB(N5697),
    .SEL(roundsel[2]),
    .O(CHOICE259)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<16>11  (
    .IA(N5698),
    .IB(N5699),
    .SEL(\c1/X[13] ),
    .O(cipherout2[17])
  );
  X_MUX2 \key2<42>110_SW01  (
    .IA(N5700),
    .IB(N5701),
    .SEL(roundsel[2]),
    .O(N5125)
  );
  X_MUX2 \key2<40>90_SW01  (
    .IA(N5702),
    .IB(N5703),
    .SEL(roundsel_2_5),
    .O(N5109)
  );
  X_MUX2 \key2<21>471  (
    .IA(N5704),
    .IB(N5705),
    .SEL(roundsel_1_6),
    .O(CHOICE980)
  );
  X_MUX2 \key2<24>1181  (
    .IA(N5706),
    .IB(N5707),
    .SEL(roundsel[3]),
    .O(CHOICE431)
  );
  X_MUX2 \key2<48>961  (
    .IA(N5708),
    .IB(N5709),
    .SEL(roundsel[2]),
    .O(CHOICE367)
  );
  X_MUX2 \key2<36>1181  (
    .IA(N5710),
    .IB(N5711),
    .SEL(roundsel[3]),
    .O(CHOICE399)
  );
  X_MUX2 \key2<23>1181  (
    .IA(N5712),
    .IB(N5713),
    .SEL(roundsel_3_3),
    .O(CHOICE908)
  );
  X_MUX2 \key2<48>110_SW01  (
    .IA(N5714),
    .IB(N5715),
    .SEL(roundsel[2]),
    .O(N5159)
  );
  X_MUX2 \c1/Mxor_X_Result<0>11  (
    .IA(N5716),
    .IB(N5717),
    .SEL(roundsel[4]),
    .O(\c1/X[1] )
  );
  X_MUX2 \key2<1>271  (
    .IA(N5718),
    .IB(N5719),
    .SEL(roundsel[1]),
    .O(CHOICE1086)
  );
  X_MUX2 \key2<44>961  (
    .IA(N5720),
    .IB(N5721),
    .SEL(roundsel_2_8),
    .O(CHOICE1789)
  );
  X_MUX2 \key2<18>110_SW01  (
    .IA(N5722),
    .IB(N5723),
    .SEL(roundsel[2]),
    .O(N5179)
  );
  X_MUX2 \key2<36>133_SW01  (
    .IA(N5724),
    .IB(N5725),
    .SEL(roundsel[3]),
    .O(N5157)
  );
  X_MUX2 \key2<16>271  (
    .IA(N5726),
    .IB(N5727),
    .SEL(roundsel_1_6),
    .O(CHOICE503)
  );
  X_MUX2 \c1/Mxor_X_Result<25>11  (
    .IA(N5728),
    .IB(N5729),
    .SEL(roundsel[4]),
    .O(\c1/X[26] )
  );
  X_MUX2 \key2<14>1181  (
    .IA(N5730),
    .IB(N5731),
    .SEL(roundsel_2_5),
    .O(CHOICE579)
  );
  X_MUX2 \key2<12>761  (
    .IA(N5732),
    .IB(N5733),
    .SEL(roundsel[2]),
    .O(CHOICE283)
  );
  X_MUX2 \key2<8>61  (
    .IA(N5734),
    .IB(N5735),
    .SEL(roundsel_2_7),
    .O(CHOICE1628)
  );
  X_MUX2 \key2<13>961  (
    .IA(N5736),
    .IB(N5737),
    .SEL(roundsel[2]),
    .O(CHOICE491)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<2>11  (
    .IA(N5738),
    .IB(N5739),
    .SEL(\c1/X[13] ),
    .O(cipherout2[3])
  );
  X_MUX2 \key2<9>471  (
    .IA(N5740),
    .IB(N5741),
    .SEL(roundsel_1_10),
    .O(CHOICE1421)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<1>11  (
    .IA(N5742),
    .IB(N5743),
    .SEL(\c1/X[1] ),
    .O(cipherout2[2])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<9>11  (
    .IA(N5744),
    .IB(N5745),
    .SEL(\c1/X[1] ),
    .O(cipherout2[10])
  );
  X_MUX2 \key2<38>110_SW01  (
    .IA(N5746),
    .IB(N5747),
    .SEL(roundsel_2_11),
    .O(N5077)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<15>11  (
    .IA(N5748),
    .IB(N5749),
    .SEL(\c1/X[1] ),
    .O(cipherout2[16])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<8>11  (
    .IA(N5750),
    .IB(N5751),
    .SEL(\c1/X[13] ),
    .O(cipherout2[9])
  );
  X_MUX2 \key2<41>110_SW01  (
    .IA(N5752),
    .IB(N5753),
    .SEL(roundsel_2_11),
    .O(N5079)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<26>11  (
    .IA(N5754),
    .IB(N5755),
    .SEL(\c1/X[13] ),
    .O(cipherout2[27])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<29>11  (
    .IA(N5756),
    .IB(N5757),
    .SEL(\c1/X[25] ),
    .O(cipherout2[30])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<22>11  (
    .IA(N5758),
    .IB(N5759),
    .SEL(\c1/X[19] ),
    .O(cipherout2[23])
  );
  X_MUX2 \_n0012<1>1051  (
    .IA(N5760),
    .IB(N5761),
    .SEL(_n0025),
    .O(N5009)
  );
  defparam \_n0012<1>1051_F .INIT = 8'h08;
  X_LUT3 \_n0012<1>1051_F  (
    .ADR0(rst_IBUF),
    .ADR1(roundsel[2]),
    .ADR2(state_FFd7),
    .O(N5760)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<12>11  (
    .IA(N5762),
    .IB(N5763),
    .SEL(\c1/X[19] ),
    .O(cipherout2[13])
  );
  X_MUX2 \key2<12>90_SW0  (
    .IA(N5764),
    .IB(N5765),
    .SEL(roundsel[3]),
    .O(N5171)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<6>11  (
    .IA(N5766),
    .IB(N5767),
    .SEL(\c1/X[19] ),
    .O(cipherout2[7])
  );
  X_MUX2 \key2<46>471  (
    .IA(N5768),
    .IB(N5769),
    .SEL(roundsel_12),
    .O(CHOICE1897)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<27>11  (
    .IA(N5770),
    .IB(N5771),
    .SEL(\c1/X[43] ),
    .O(cipherout2[28])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<11>11  (
    .IA(N5772),
    .IB(N5773),
    .SEL(\c1/X[43] ),
    .O(cipherout2[12])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<23>11  (
    .IA(N5774),
    .IB(N5775),
    .SEL(\c1/X[1] ),
    .O(cipherout2[24])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<10>11  (
    .IA(N5776),
    .IB(N5777),
    .SEL(\c1/X[37] ),
    .O(cipherout2[11])
  );
  X_MUX2 \key2<8>271  (
    .IA(N5778),
    .IB(N5779),
    .SEL(roundsel_1_10),
    .O(CHOICE1621)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<5>11  (
    .IA(N5780),
    .IB(N5781),
    .SEL(\c1/X[43] ),
    .O(cipherout2[6])
  );
  X_MUX2 \key2<40>761  (
    .IA(N5782),
    .IB(N5783),
    .SEL(roundsel_2_8),
    .O(CHOICE1705)
  );
  X_MUX2 \c1/Mxor_OUTR_Result<18>11  (
    .IA(N5784),
    .IB(N5785),
    .SEL(\c1/X[25] ),
    .O(cipherout2[19])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<0>11  (
    .IA(N5786),
    .IB(N5787),
    .SEL(\c1/X[37] ),
    .O(cipherout2[1])
  );
  X_MUX2 \c1/Mxor_OUTR_Result<17>11  (
    .IA(N5788),
    .IB(N5789),
    .SEL(\c1/X[43] ),
    .O(cipherout2[18])
  );
  X_MUX2 \key2<2>961  (
    .IA(N5790),
    .IB(N5791),
    .SEL(roundsel_2_8),
    .O(CHOICE1733)
  );
  X_MUX2 \key2<26>271  (
    .IA(N5792),
    .IB(N5793),
    .SEL(roundsel_1_6),
    .O(CHOICE1645)
  );
  X_MUX2 \key2<29>1181  (
    .IA(N5794),
    .IB(N5795),
    .SEL(roundsel_2_8),
    .O(CHOICE1553)
  );
  X_MUX2 \key2<15>1191  (
    .IA(N5796),
    .IB(N5797),
    .SEL(roundsel_3_14),
    .O(CHOICE611)
  );
  X_MUX2 \key2<20>961  (
    .IA(N5798),
    .IB(N5799),
    .SEL(roundsel_2_12),
    .O(CHOICE964)
  );
  X_MUX2 \key2<37>271  (
    .IA(N5800),
    .IB(N5801),
    .SEL(roundsel[1]),
    .O(CHOICE1162)
  );
  X_MUX2 \key2<11>110_SW01  (
    .IA(N5802),
    .IB(N5803),
    .SEL(roundsel_2_13),
    .O(N5061)
  );
  X_MUX2 \key2<25>271  (
    .IA(N5804),
    .IB(N5805),
    .SEL(roundsel_1_6),
    .O(CHOICE1134)
  );
  X_MUX2 \key2<11>961  (
    .IA(N5806),
    .IB(N5807),
    .SEL(roundsel_2_13),
    .O(CHOICE1521)
  );
  X_MUX2 \key2<39>90_SW01  (
    .IA(N5808),
    .IB(N5809),
    .SEL(roundsel_2_11),
    .O(N5107)
  );
  X_MUX2 \key2<23>133_SW01  (
    .IA(N5810),
    .IB(N5811),
    .SEL(roundsel_33),
    .O(N5069)
  );
  X_MUX2 \key2<30>133_SW01  (
    .IA(N5812),
    .IB(N5813),
    .SEL(roundsel[2]),
    .O(N5155)
  );
  X_MUX2 \key2<46>1191  (
    .IA(N5814),
    .IB(N5815),
    .SEL(roundsel_2_12),
    .O(CHOICE1913)
  );
  X_MUX2 \key2<13>271  (
    .IA(N5816),
    .IB(N5817),
    .SEL(roundsel[1]),
    .O(CHOICE475)
  );
  X_MUX2 \key2<42>961  (
    .IA(N5818),
    .IB(N5819),
    .SEL(roundsel[2]),
    .O(CHOICE311)
  );
  X_MUX2 \key2<10>961  (
    .IA(N5820),
    .IB(N5821),
    .SEL(roundsel_2_13),
    .O(CHOICE1262)
  );
  X_MUX2 \key2<15>471  (
    .IA(N5822),
    .IB(N5823),
    .SEL(roundsel_1_22),
    .O(CHOICE595)
  );
  X_MUX2 \key2<9>1191  (
    .IA(N5824),
    .IB(N5825),
    .SEL(roundsel_2_12),
    .O(CHOICE1437)
  );
  X_MUX2 \key2<27>471  (
    .IA(N5826),
    .IB(N5827),
    .SEL(roundsel_1_22),
    .O(CHOICE1320)
  );
  X_MUX2 \c1/Mxor_X_Result<31>11  (
    .IA(N5828),
    .IB(N5829),
    .SEL(roundsel_43),
    .O(\c1/X[32] )
  );
  X_MUX2 \key2<24>133_SW01  (
    .IA(N5830),
    .IB(N5831),
    .SEL(roundsel[3]),
    .O(N5123)
  );
  X_MUX2 \key2<27>1411  (
    .IA(N5832),
    .IB(N5833),
    .SEL(roundsel_2_8),
    .O(CHOICE1340)
  );
  X_MUX2 \key2<10>110_SW01  (
    .IA(N5834),
    .IB(N5835),
    .SEL(roundsel_2_13),
    .O(N5059)
  );
  X_MUX2 \key2<2>110_SW01  (
    .IA(N5836),
    .IB(N5837),
    .SEL(roundsel_2_5),
    .O(N5087)
  );
  X_MUX2 \key2<5>110_SW01  (
    .IA(N5838),
    .IB(N5839),
    .SEL(roundsel_3_15),
    .O(N5091)
  );
  X_MUX2 \key2<7>761  (
    .IA(N5840),
    .IB(N5841),
    .SEL(roundsel_2_13),
    .O(CHOICE1074)
  );
  X_MUX2 \key2<33>110_SW01  (
    .IA(N5842),
    .IB(N5843),
    .SEL(roundsel_2_4),
    .O(N5073)
  );
  X_MUX2 \key2<45>1191  (
    .IA(N5844),
    .IB(N5845),
    .SEL(roundsel_4_7),
    .O(CHOICE1881)
  );
  X_MUX2 \key2<5>961  (
    .IA(N5846),
    .IB(N5847),
    .SEL(roundsel_3_15),
    .O(CHOICE1405)
  );
  X_MUX2 \key2<14>133_SW01  (
    .IA(N5848),
    .IB(N5849),
    .SEL(roundsel_2_11),
    .O(N5063)
  );
  X_MUX2 \key2<43>271  (
    .IA(N5850),
    .IB(N5851),
    .SEL(roundsel[1]),
    .O(CHOICE1190)
  );
  X_MUX2 \c1/Mxor_X_Result<15>11  (
    .IA(N5852),
    .IB(N5853),
    .SEL(roundsel[4]),
    .O(\c1/X[16] )
  );
  X_MUX2 \key2<28>471  (
    .IA(N5854),
    .IB(N5855),
    .SEL(roundsel_1_22),
    .O(CHOICE1833)
  );
  X_MUX2 \key2<17>1191  (
    .IA(N5856),
    .IB(N5857),
    .SEL(roundsel_33),
    .O(CHOICE547)
  );
  X_MUX2 \key2<20>110_SW01  (
    .IA(N5858),
    .IB(N5859),
    .SEL(roundsel_2_12),
    .O(N5065)
  );
  X_MUX2 \c1/u4/Mrom_dout_inst_mux_f5_291  (
    .IA(N5860),
    .IB(N5861),
    .SEL(\c1/X[25] ),
    .O(\c1/u4/Mrom_dout_N7 )
  );
  X_MUX2 \c1/u4/Mrom_dout_inst_mux_f5_281  (
    .IA(N5862),
    .IB(N5863),
    .SEL(\c1/X[25] ),
    .O(\c1/u4/Mrom_dout_N6 )
  );
  X_MUX2 \roundsel<2>_mmx_out331  (
    .IA(N5864),
    .IB(N5865),
    .SEL(roundsel[2]),
    .O(\MUX_BLOCK_roundsel<2>_mmx_out33 )
  );
  X_MUX2 \c1/u4/Mrom_dout_inst_mux_f5_251  (
    .IA(N5866),
    .IB(N5867),
    .SEL(\c1/X[25] ),
    .O(\c1/u4/Mrom_dout_N1 )
  );
  X_MUX2 \c1/u4/Mrom_dout_inst_mux_f5_241  (
    .IA(N5868),
    .IB(N5869),
    .SEL(\c1/X[25] ),
    .O(\c1/u4/Mrom_dout_N0 )
  );
  X_MUX2 \c1/u6/Mrom_dout_inst_mux_f5_111  (
    .IA(N5870),
    .IB(N5871),
    .SEL(\c1/X[37] ),
    .O(\c1/u6/Mrom_dout_N4 )
  );
  X_MUX2 \c1/u6/Mrom_dout_inst_mux_f5_101  (
    .IA(N5872),
    .IB(N5873),
    .SEL(\c1/X[37] ),
    .O(\c1/u6/Mrom_dout_N3 )
  );
  X_MUX2 \c1/Mxor_OUTR_Result<25>11  (
    .IA(N5874),
    .IB(N5875),
    .SEL(\c1/X[37] ),
    .O(cipherout2[26])
  );
  X_MUX2 \roundsel<2>_mmx_out241  (
    .IA(N5876),
    .IB(N5877),
    .SEL(roundsel_2_7),
    .O(\MUX_BLOCK_roundsel<2>_mmx_out24 )
  );
  X_MUX2 \key2<31>15  (
    .IA(N5878),
    .IB(N5879),
    .SEL(roundsel_2_10),
    .O(CHOICE1106)
  );
  X_MUX2 \key2<26>12  (
    .IA(N5880),
    .IB(N5881),
    .SEL(roundsel_3_11),
    .O(CHOICE1639)
  );
  X_MUX2 \key2<8>12  (
    .IA(N5882),
    .IB(N5883),
    .SEL(roundsel_3_13),
    .O(CHOICE1615)
  );
  X_MUX2 \key2<37>12_SW0  (
    .IA(N5884),
    .IB(N5885),
    .SEL(roundsel_3_6),
    .O(N5175)
  );
  X_MUX2 \key2<43>12_SW0  (
    .IA(N5886),
    .IB(N5887),
    .SEL(roundsel_3_6),
    .O(N5177)
  );
  X_MUX2 \key2<13>12_SW0  (
    .IA(N5888),
    .IB(N5889),
    .SEL(roundsel_3_6),
    .O(N5195)
  );
  X_MUX2 \key2<7>15  (
    .IA(N5890),
    .IB(N5891),
    .SEL(roundsel_2_10),
    .O(CHOICE1058)
  );
  X_MUX2 \key2<26>61  (
    .IA(N5892),
    .IB(N5893),
    .SEL(roundsel_23),
    .O(CHOICE1652)
  );
  X_MUX2 \key2<31>12  (
    .IA(N5894),
    .IB(N5895),
    .SEL(roundsel_2_10),
    .O(CHOICE1104)
  );
  X_MUX2 \key2<7>12  (
    .IA(N5896),
    .IB(N5897),
    .SEL(roundsel_24),
    .O(CHOICE1056)
  );
  X_OPAD \dataout<1>  (
    .PAD(dataout[1])
  );
  X_IPAD \key<52>  (
    .PAD(key[52])
  );
  X_IPAD \datain<6>  (
    .PAD(datain[6])
  );
  X_IPAD \datain<26>  (
    .PAD(datain[26])
  );
  X_OPAD \dataout<23>  (
    .PAD(dataout[23])
  );
  X_IPAD \key<36>  (
    .PAD(key[36])
  );
  X_IPAD \datain<58>  (
    .PAD(datain[58])
  );
  X_IPAD \datain<2>  (
    .PAD(datain[2])
  );
  X_IPAD \datain<4>  (
    .PAD(datain[4])
  );
  X_IPAD \datain<60>  (
    .PAD(datain[60])
  );
  X_IPAD \key<60>  (
    .PAD(key[60])
  );
  X_OPAD \dataout<4>  (
    .PAD(dataout[4])
  );
  X_OPAD \dataout<48>  (
    .PAD(dataout[48])
  );
  X_OPAD \dataout<43>  (
    .PAD(dataout[43])
  );
  X_IPAD \key<8>  (
    .PAD(key[8])
  );
  X_OPAD \dataout<25>  (
    .PAD(dataout[25])
  );
  X_OPAD \dataout<49>  (
    .PAD(dataout[49])
  );
  X_IPAD \key<62>  (
    .PAD(key[62])
  );
  X_OPAD \dataout<31>  (
    .PAD(dataout[31])
  );
  X_OPAD \dataout<24>  (
    .PAD(dataout[24])
  );
  X_IPAD \key<64>  (
    .PAD(key[64])
  );
  X_OPAD \dataout<35>  (
    .PAD(dataout[35])
  );
  X_OPAD \dataout<33>  (
    .PAD(dataout[33])
  );
  X_OPAD \dataout<46>  (
    .PAD(dataout[46])
  );
  X_IPAD \datain<23>  (
    .PAD(datain[23])
  );
  X_OPAD \dataout<26>  (
    .PAD(dataout[26])
  );
  X_OPAD \dataout<17>  (
    .PAD(dataout[17])
  );
  X_IPAD \key<63>  (
    .PAD(key[63])
  );
  X_OPAD \dataout<45>  (
    .PAD(dataout[45])
  );
  X_OPAD \dataout<40>  (
    .PAD(dataout[40])
  );
  X_OPAD \dataout<42>  (
    .PAD(dataout[42])
  );
  X_OPAD \dataout<6>  (
    .PAD(dataout[6])
  );
  X_OPAD \dataout<3>  (
    .PAD(dataout[3])
  );
  X_OPAD \dataout<51>  (
    .PAD(dataout[51])
  );
  X_IPAD \datain<19>  (
    .PAD(datain[19])
  );
  X_IPAD \key<61>  (
    .PAD(key[61])
  );
  X_OPAD \dataout<28>  (
    .PAD(dataout[28])
  );
  X_OPAD \dataout<5>  (
    .PAD(dataout[5])
  );
  X_OPAD \dataout<37>  (
    .PAD(dataout[37])
  );
  X_OPAD \dataout<36>  (
    .PAD(dataout[36])
  );
  X_OPAD \dataout<30>  (
    .PAD(dataout[30])
  );
  X_OPAD \dataout<39>  (
    .PAD(dataout[39])
  );
  X_OPAD \dataout<32>  (
    .PAD(dataout[32])
  );
  X_OPAD \dataout<29>  (
    .PAD(dataout[29])
  );
  X_OPAD \dataout<27>  (
    .PAD(dataout[27])
  );
  X_OPAD \dataout<34>  (
    .PAD(dataout[34])
  );
  X_OPAD \dataout<47>  (
    .PAD(dataout[47])
  );
  X_OPAD \dataout<38>  (
    .PAD(dataout[38])
  );
  X_IPAD \datain<55>  (
    .PAD(datain[55])
  );
  X_IPAD \key<20>  (
    .PAD(key[20])
  );
  X_OPAD \dataout<41>  (
    .PAD(dataout[41])
  );
  X_OPAD \dataout<50>  (
    .PAD(dataout[50])
  );
  X_OPAD \dataout<44>  (
    .PAD(dataout[44])
  );
  X_IPAD \key<55>  (
    .PAD(key[55])
  );
  X_IPAD \datain<36>  (
    .PAD(datain[36])
  );
  X_IPAD \datain<56>  (
    .PAD(datain[56])
  );
  X_IPAD \datain<42>  (
    .PAD(datain[42])
  );
  X_IPAD \datain<13>  (
    .PAD(datain[13])
  );
  X_IPAD \key<5>  (
    .PAD(key[5])
  );
  X_IPAD rst_248 (
    .PAD(rst)
  );
  X_IPAD \key<23>  (
    .PAD(key[23])
  );
  X_OPAD \dataout<2>  (
    .PAD(dataout[2])
  );
  X_OPAD \ready.PAD  (
    .PAD(ready)
  );
  X_IPAD \datain<34>  (
    .PAD(datain[34])
  );
  X_IPAD \key<21>  (
    .PAD(key[21])
  );
  X_IPAD \datain<57>  (
    .PAD(datain[57])
  );
  X_OPAD \dataout<15>  (
    .PAD(dataout[15])
  );
  X_IPAD \datain<39>  (
    .PAD(datain[39])
  );
  X_IPAD \key<31>  (
    .PAD(key[31])
  );
  X_IPAD \datain<11>  (
    .PAD(datain[11])
  );
  X_IPAD \key<19>  (
    .PAD(key[19])
  );
  X_IPAD \datain<9>  (
    .PAD(datain[9])
  );
  X_OPAD \dataout<11>  (
    .PAD(dataout[11])
  );
  X_OPAD \dataout<14>  (
    .PAD(dataout[14])
  );
  X_IPAD \datain<7>  (
    .PAD(datain[7])
  );
  X_IPAD \datain<8>  (
    .PAD(datain[8])
  );
  X_OPAD \dataout<61>  (
    .PAD(dataout[61])
  );
  X_OPAD \dataout<7>  (
    .PAD(dataout[7])
  );
  X_IPAD \key<32>  (
    .PAD(key[32])
  );
  X_IPAD \datain<50>  (
    .PAD(datain[50])
  );
  X_OPAD \dataout<63>  (
    .PAD(dataout[63])
  );
  X_IPAD \key<39>  (
    .PAD(key[39])
  );
  X_IPAD \datain<5>  (
    .PAD(datain[5])
  );
  X_IPAD \datain<30>  (
    .PAD(datain[30])
  );
  X_IPAD \datain<47>  (
    .PAD(datain[47])
  );
  X_IPAD \datain<49>  (
    .PAD(datain[49])
  );
  X_OPAD \dataout<64>  (
    .PAD(dataout[64])
  );
  X_IPAD \datain<59>  (
    .PAD(datain[59])
  );
  X_IPAD \datain<48>  (
    .PAD(datain[48])
  );
  X_IPAD \key<13>  (
    .PAD(key[13])
  );
  X_OPAD \dataout<8>  (
    .PAD(dataout[8])
  );
  X_IPAD \key<47>  (
    .PAD(key[47])
  );
  X_OPAD \dataout<52>  (
    .PAD(dataout[52])
  );
  X_IPAD \key<29>  (
    .PAD(key[29])
  );
  X_IPAD clk_249 (
    .PAD(clk)
  );
  X_IPAD \datain<29>  (
    .PAD(datain[29])
  );
  X_IPAD \key<3>  (
    .PAD(key[3])
  );
  X_OPAD \dataout<9>  (
    .PAD(dataout[9])
  );
  X_IPAD \datain<35>  (
    .PAD(datain[35])
  );
  X_IPAD \datain<28>  (
    .PAD(datain[28])
  );
  X_IPAD \datain<1>  (
    .PAD(datain[1])
  );
  X_IPAD \key<6>  (
    .PAD(key[6])
  );
  X_IPAD \key<53>  (
    .PAD(key[53])
  );
  X_IPAD \datain<44>  (
    .PAD(datain[44])
  );
  X_OPAD \dataout<56>  (
    .PAD(dataout[56])
  );
  X_OPAD \dataout<21>  (
    .PAD(dataout[21])
  );
  X_OPAD \dataout<62>  (
    .PAD(dataout[62])
  );
  X_OPAD \dataout<57>  (
    .PAD(dataout[57])
  );
  X_OPAD \dataout<19>  (
    .PAD(dataout[19])
  );
  X_OPAD \dataout<60>  (
    .PAD(dataout[60])
  );
  X_IPAD \key<18>  (
    .PAD(key[18])
  );
  X_OPAD \dataout<58>  (
    .PAD(dataout[58])
  );
  X_IPAD \datain<63>  (
    .PAD(datain[63])
  );
  X_IPAD \key<30>  (
    .PAD(key[30])
  );
  X_IPAD \datain<64>  (
    .PAD(datain[64])
  );
  X_IPAD \key<34>  (
    .PAD(key[34])
  );
  X_IPAD \datain<20>  (
    .PAD(datain[20])
  );
  X_OPAD \dataout<10>  (
    .PAD(dataout[10])
  );
  X_IPAD \key<50>  (
    .PAD(key[50])
  );
  X_IPAD \key<42>  (
    .PAD(key[42])
  );
  X_IPAD \key<2>  (
    .PAD(key[2])
  );
  X_IPAD \key<35>  (
    .PAD(key[35])
  );
  X_IPAD \key<26>  (
    .PAD(key[26])
  );
  X_OPAD \dataout<55>  (
    .PAD(dataout[55])
  );
  X_IPAD \datain<53>  (
    .PAD(datain[53])
  );
  X_IPAD \datain<25>  (
    .PAD(datain[25])
  );
  X_IPAD \key<16>  (
    .PAD(key[16])
  );
  X_IPAD \datain<37>  (
    .PAD(datain[37])
  );
  X_IPAD \key<40>  (
    .PAD(key[40])
  );
  X_IPAD \key<37>  (
    .PAD(key[37])
  );
  X_IPAD \datain<51>  (
    .PAD(datain[51])
  );
  X_IPAD \datain<22>  (
    .PAD(datain[22])
  );
  X_IPAD \key<24>  (
    .PAD(key[24])
  );
  X_IPAD \key<54>  (
    .PAD(key[54])
  );
  X_IPAD \datain<14>  (
    .PAD(datain[14])
  );
  X_IPAD \datain<33>  (
    .PAD(datain[33])
  );
  X_OPAD \dataout<54>  (
    .PAD(dataout[54])
  );
  X_IPAD \datain<17>  (
    .PAD(datain[17])
  );
  X_IPAD \datain<46>  (
    .PAD(datain[46])
  );
  X_IPAD \key<7>  (
    .PAD(key[7])
  );
  X_IPAD \datain<38>  (
    .PAD(datain[38])
  );
  X_OPAD \dataout<12>  (
    .PAD(dataout[12])
  );
  X_OPAD \dataout<22>  (
    .PAD(dataout[22])
  );
  X_IPAD \datain<62>  (
    .PAD(datain[62])
  );
  X_IPAD \datain<3>  (
    .PAD(datain[3])
  );
  X_IPAD \datain<15>  (
    .PAD(datain[15])
  );
  X_IPAD \key<28>  (
    .PAD(key[28])
  );
  X_IPAD \datain<12>  (
    .PAD(datain[12])
  );
  X_IPAD \datain<16>  (
    .PAD(datain[16])
  );
  X_IPAD \key<56>  (
    .PAD(key[56])
  );
  X_IPAD \key<46>  (
    .PAD(key[46])
  );
  X_IPAD \datain<18>  (
    .PAD(datain[18])
  );
  X_IPAD \datain<43>  (
    .PAD(datain[43])
  );
  X_IPAD \datain<41>  (
    .PAD(datain[41])
  );
  X_OPAD \dataout<16>  (
    .PAD(dataout[16])
  );
  X_IPAD \key<58>  (
    .PAD(key[58])
  );
  X_IPAD \datain<54>  (
    .PAD(datain[54])
  );
  X_IPAD \key<51>  (
    .PAD(key[51])
  );
  X_IPAD \key<22>  (
    .PAD(key[22])
  );
  X_OPAD \dataout<59>  (
    .PAD(dataout[59])
  );
  X_IPAD \datain<10>  (
    .PAD(datain[10])
  );
  X_OPAD \dataout<13>  (
    .PAD(dataout[13])
  );
  X_IPAD \datain<32>  (
    .PAD(datain[32])
  );
  X_IPAD \key<11>  (
    .PAD(key[11])
  );
  X_OPAD \dataout<18>  (
    .PAD(dataout[18])
  );
  X_IPAD \key<43>  (
    .PAD(key[43])
  );
  X_IPAD \datain<40>  (
    .PAD(datain[40])
  );
  X_IPAD \key<38>  (
    .PAD(key[38])
  );
  X_IPAD \datain<45>  (
    .PAD(datain[45])
  );
  X_IPAD \datain<24>  (
    .PAD(datain[24])
  );
  X_IPAD \datain<31>  (
    .PAD(datain[31])
  );
  X_IPAD \key<4>  (
    .PAD(key[4])
  );
  X_IPAD \datain<61>  (
    .PAD(datain[61])
  );
  X_IPAD \datain<21>  (
    .PAD(datain[21])
  );
  X_IPAD \key<48>  (
    .PAD(key[48])
  );
  X_OPAD \dataout<53>  (
    .PAD(dataout[53])
  );
  X_IPAD \datain<52>  (
    .PAD(datain[52])
  );
  X_IPAD \key<59>  (
    .PAD(key[59])
  );
  X_IPAD flag_250 (
    .PAD(flag)
  );
  X_IPAD \key<27>  (
    .PAD(key[27])
  );
  X_IPAD \key<45>  (
    .PAD(key[45])
  );
  X_IPAD \key<14>  (
    .PAD(key[14])
  );
  X_IPAD \key<15>  (
    .PAD(key[15])
  );
  X_IPAD \datain<27>  (
    .PAD(datain[27])
  );
  X_IPAD \key<12>  (
    .PAD(key[12])
  );
  X_IPAD \key<44>  (
    .PAD(key[44])
  );
  X_OPAD \dataout<20>  (
    .PAD(dataout[20])
  );
  X_IPAD \key<10>  (
    .PAD(key[10])
  );
  X_BUF \key2<7>90/LUT4_D_BUF  (
    .I(\key2[7] ),
    .O(N5898)
  );
  defparam \key2<7>90 .INIT = 16'hFAF8;
  X_LUT4 \key2<7>90  (
    .ADR0(roundsel[4]),
    .ADR1(CHOICE1056),
    .ADR2(CHOICE1074),
    .ADR3(CHOICE1058),
    .O(\key2[7] )
  );
  X_BUF \key2<7>12_F/LUT4_L_BUF  (
    .I(\key2<7>12_F/O ),
    .O(N5896)
  );
  defparam \key2<7>12_F .INIT = 16'hA280;
  X_LUT4 \key2<7>12_F  (
    .ADR0(roundsel_3_6),
    .ADR1(roundsel_1_18),
    .ADR2(\key1[44] ),
    .ADR3(\key1[28] ),
    .O(\key2<7>12_F/O )
  );
  X_BUF \_n0013<6>22/LUT4_L_BUF  (
    .I(\_n0013<6>22/O ),
    .O(_n0013[6])
  );
  defparam \_n0013<6>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<6>22  (
    .ADR0(CHOICE633),
    .ADR1(N5450),
    .ADR2(cipherout2[7]),
    .ADR3(_n0025),
    .O(\_n0013<6>22/O )
  );
  X_BUF \key2<22>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<22>110_SW01_G/O ),
    .O(N5621)
  );
  defparam \key2<22>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<22>110_SW01_G  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out42 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out39 ),
    .O(\key2<22>110_SW01_G/O )
  );
  X_BUF \_n0013<8>22/LUT4_L_BUF  (
    .I(\_n0013<8>22/O ),
    .O(_n0013[8])
  );
  defparam \_n0013<8>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<8>22  (
    .ADR0(CHOICE642),
    .ADR1(N5452),
    .ADR2(cipherout2[9]),
    .ADR3(_n0025),
    .O(\_n0013<8>22/O )
  );
  X_BUF \_n0013<13>20/LUT4_L_BUF  (
    .I(\_n0013<13>20/O ),
    .O(_n0013[13])
  );
  defparam \_n0013<13>20 .INIT = 16'hFFEA;
  X_LUT4 \_n0013<13>20  (
    .ADR0(CHOICE2017),
    .ADR1(_n0025),
    .ADR2(cipherout2[14]),
    .ADR3(N5432),
    .O(\_n0013<13>20/O )
  );
  X_BUF \_n0013<10>22/LUT4_L_BUF  (
    .I(\_n0013<10>22/O ),
    .O(_n0013[10])
  );
  defparam \_n0013<10>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<10>22  (
    .ADR0(CHOICE651),
    .ADR1(N5454),
    .ADR2(cipherout2[11]),
    .ADR3(_n0025),
    .O(\_n0013<10>22/O )
  );
  X_BUF \key2<4>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<4>110_SW01_G/O ),
    .O(N5623)
  );
  defparam \key2<4>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<4>110_SW01_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out68 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out44 ),
    .O(\key2<4>110_SW01_G/O )
  );
  X_BUF \_n0013<0>22/LUT4_L_BUF  (
    .I(\_n0013<0>22/O ),
    .O(_n0013[0])
  );
  defparam \_n0013<0>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<0>22  (
    .ADR0(CHOICE660),
    .ADR1(N5456),
    .ADR2(cipherout2[1]),
    .ADR3(_n0025),
    .O(\_n0013<0>22/O )
  );
  X_BUF \_n0013<2>22/LUT4_L_BUF  (
    .I(\_n0013<2>22/O ),
    .O(_n0013[2])
  );
  defparam \_n0013<2>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<2>22  (
    .ADR0(CHOICE669),
    .ADR1(N5458),
    .ADR2(cipherout2[3]),
    .ADR3(_n0025),
    .O(\_n0013<2>22/O )
  );
  X_BUF \_n0013<7>20/LUT4_L_BUF  (
    .I(\_n0013<7>20/O ),
    .O(_n0013[7])
  );
  defparam \_n0013<7>20 .INIT = 16'hFFEA;
  X_LUT4 \_n0013<7>20  (
    .ADR0(CHOICE1918),
    .ADR1(\state_FFd3-In ),
    .ADR2(cipherout2[1]),
    .ADR3(N5430),
    .O(\_n0013<7>20/O )
  );
  X_BUF \_n0013<4>22/LUT4_L_BUF  (
    .I(\_n0013<4>22/O ),
    .O(_n0013[4])
  );
  defparam \_n0013<4>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<4>22  (
    .ADR0(CHOICE675),
    .ADR1(CHOICE680),
    .ADR2(N5910),
    .ADR3(_n0025),
    .O(\_n0013<4>22/O )
  );
  X_BUF \key2<3>1181_G/LUT4_L_BUF  (
    .I(\key2<3>1181_G/O ),
    .O(N5625)
  );
  defparam \key2<3>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<3>1181_G  (
    .ADR0(roundsel_4_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out60 ),
    .ADR2(roundsel_2_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out49 ),
    .O(\key2<3>1181_G/O )
  );
  X_BUF \_n0013<63>22/LUT4_L_BUF  (
    .I(\_n0013<63>22/O ),
    .O(_n0013[63])
  );
  defparam \_n0013<63>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<63>22  (
    .ADR0(CHOICE686),
    .ADR1(N5460),
    .ADR2(N5907),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<63>22/O )
  );
  X_BUF \_n0013<32>21/LUT3_L_BUF  (
    .I(\_n0013<32>21/O ),
    .O(_n0013[32])
  );
  defparam \_n0013<32>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<32>21  (
    .ADR0(CHOICE149),
    .ADR1(data1[33]),
    .ADR2(N01),
    .O(\_n0013<32>21/O )
  );
  X_BUF \_n0013<61>22/LUT4_L_BUF  (
    .I(\_n0013<61>22/O ),
    .O(_n0013[61])
  );
  defparam \_n0013<61>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<61>22  (
    .ADR0(CHOICE695),
    .ADR1(N5462),
    .ADR2(cipherout2[16]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<61>22/O )
  );
  X_BUF \key2<32>271_G/LUT4_L_BUF  (
    .I(\key2<32>271_G/O ),
    .O(N5627)
  );
  defparam \key2<32>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<32>271_G  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[55] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[54] ),
    .O(\key2<32>271_G/O )
  );
  X_BUF \_n0013<59>22/LUT4_L_BUF  (
    .I(\_n0013<59>22/O ),
    .O(_n0013[59])
  );
  defparam \_n0013<59>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<59>22  (
    .ADR0(CHOICE704),
    .ADR1(N5464),
    .ADR2(cipherout2[24]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<59>22/O )
  );
  X_BUF \_n0013<48>5/LUT4_L_BUF  (
    .I(\_n0013<48>5/O ),
    .O(CHOICE91)
  );
  defparam \_n0013<48>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<48>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[4]),
    .ADR2(state_FFd8),
    .ADR3(datain_49_IBUF),
    .O(\_n0013<48>5/O )
  );
  X_BUF \_n0013<57>22/LUT4_L_BUF  (
    .I(\_n0013<57>22/O ),
    .O(_n0013[57])
  );
  defparam \_n0013<57>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<57>22  (
    .ADR0(CHOICE713),
    .ADR1(N5440),
    .ADR2(cipherout2[32]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<57>22/O )
  );
  X_BUF \_n0013<55>22/LUT4_L_BUF  (
    .I(\_n0013<55>22/O ),
    .O(_n0013[55])
  );
  defparam \_n0013<55>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<55>22  (
    .ADR0(CHOICE722),
    .ADR1(N5466),
    .ADR2(cipherout2[7]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<55>22/O )
  );
  X_BUF \_n0013<53>22/LUT4_L_BUF  (
    .I(\_n0013<53>22/O ),
    .O(_n0013[53])
  );
  defparam \_n0013<53>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<53>22  (
    .ADR0(CHOICE733),
    .ADR1(CHOICE734),
    .ADR2(N5909),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<53>22/O )
  );
  X_BUF \_n0013<57>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<57>22_SW0/O ),
    .O(N5440)
  );
  defparam \_n0013<57>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<57>22_SW0  (
    .ADR0(data1[26]),
    .ADR1(_n0025),
    .ADR2(data1[58]),
    .ADR3(N01),
    .O(\_n0013<57>22_SW0/O )
  );
  X_BUF \_n0013<51>22/LUT4_L_BUF  (
    .I(\_n0013<51>22/O ),
    .O(_n0013[51])
  );
  defparam \_n0013<51>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<51>22  (
    .ADR0(CHOICE740),
    .ADR1(N5468),
    .ADR2(cipherout2[23]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<51>22/O )
  );
  X_BUF \_n0013<8>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<8>22_SW0/O ),
    .O(N5452)
  );
  defparam \_n0013<8>22_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<8>22_SW0  (
    .ADR0(data1[26]),
    .ADR1(data1[9]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<8>22_SW0/O )
  );
  X_BUF \_n0013<49>22/LUT4_L_BUF  (
    .I(\_n0013<49>22/O ),
    .O(_n0013[49])
  );
  defparam \_n0013<49>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<49>22  (
    .ADR0(CHOICE751),
    .ADR1(CHOICE752),
    .ADR2(N5915),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<49>22/O )
  );
  X_BUF \key2<47>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<47>110_SW01_G/O ),
    .O(N5629)
  );
  defparam \key2<47>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<47>110_SW01_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out82 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out80 ),
    .O(\key2<47>110_SW01_G/O )
  );
  X_BUF \_n0013<47>22/LUT4_L_BUF  (
    .I(\_n0013<47>22/O ),
    .O(_n0013[47])
  );
  defparam \_n0013<47>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<47>22  (
    .ADR0(CHOICE758),
    .ADR1(N5470),
    .ADR2(cipherout2[6]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<47>22/O )
  );
  X_BUF \_n0013<45>17/LUT4_L_BUF  (
    .I(\_n0013<45>17/O ),
    .O(_n0013[45])
  );
  defparam \_n0013<45>17 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<45>17  (
    .ADR0(CHOICE624),
    .ADR1(CHOICE626),
    .ADR2(N5908),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<45>17/O )
  );
  X_BUF \key2<28>1191_G/LUT4_L_BUF  (
    .I(\key2<28>1191_G/O ),
    .O(N5631)
  );
  defparam \key2<28>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<28>1191_G  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .ADR2(roundsel_3_15),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .O(\key2<28>1191_G/O )
  );
  X_BUF \_n0013<43>22/LUT4_L_BUF  (
    .I(\_n0013<43>22/O ),
    .O(_n0013[43])
  );
  defparam \_n0013<43>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<43>22  (
    .ADR0(CHOICE767),
    .ADR1(N5442),
    .ADR2(N5912),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<43>22/O )
  );
  X_BUF \_n0013<41>22/LUT4_L_BUF  (
    .I(\_n0013<41>22/O ),
    .O(_n0013[41])
  );
  defparam \_n0013<41>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<41>22  (
    .ADR0(CHOICE776),
    .ADR1(N5472),
    .ADR2(cipherout2[30]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<41>22/O )
  );
  X_BUF \_n0013<39>22/LUT4_L_BUF  (
    .I(\_n0013<39>22/O ),
    .O(_n0013[39])
  );
  defparam \_n0013<39>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<39>22  (
    .ADR0(CHOICE787),
    .ADR1(CHOICE788),
    .ADR2(cipherout2[5]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<39>22/O )
  );
  X_BUF \_n0013<37>22/LUT4_L_BUF  (
    .I(\_n0013<37>22/O ),
    .O(_n0013[37])
  );
  defparam \_n0013<37>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<37>22  (
    .ADR0(CHOICE794),
    .ADR1(N5474),
    .ADR2(cipherout2[13]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<37>22/O )
  );
  X_BUF \_n0013<35>22/LUT4_L_BUF  (
    .I(\_n0013<35>22/O ),
    .O(_n0013[35])
  );
  defparam \_n0013<35>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<35>22  (
    .ADR0(CHOICE803),
    .ADR1(N5476),
    .ADR2(N5911),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<35>22/O )
  );
  X_BUF \_n0013<34>5/LUT4_L_BUF  (
    .I(\_n0013<34>5/O ),
    .O(CHOICE154)
  );
  defparam \_n0013<34>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<34>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[24]),
    .ADR2(state_FFd8),
    .ADR3(datain_35_IBUF),
    .O(\_n0013<34>5/O )
  );
  X_BUF \_n0013<33>22/LUT4_L_BUF  (
    .I(\_n0013<33>22/O ),
    .O(_n0013[33])
  );
  defparam \_n0013<33>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<33>22  (
    .ADR0(CHOICE812),
    .ADR1(N5444),
    .ADR2(N5914),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<33>22/O )
  );
  X_BUF \_n0013<48>14/LUT3_L_BUF  (
    .I(\_n0013<48>14/O ),
    .O(CHOICE95)
  );
  defparam \_n0013<48>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<48>14  (
    .ADR0(CHOICE93),
    .ADR1(data1[31]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<48>14/O )
  );
  X_BUF \_n0013<30>22/LUT4_L_BUF  (
    .I(\_n0013<30>22/O ),
    .O(_n0013[30])
  );
  defparam \_n0013<30>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<30>22  (
    .ADR0(CHOICE819),
    .ADR1(CHOICE824),
    .ADR2(cipherout2[31]),
    .ADR3(_n0025),
    .O(\_n0013<30>22/O )
  );
  X_BUF \_n0013<28>22/LUT4_L_BUF  (
    .I(\_n0013<28>22/O ),
    .O(_n0013[28])
  );
  defparam \_n0013<28>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<28>22  (
    .ADR0(CHOICE831),
    .ADR1(N5446),
    .ADR2(cipherout2[29]),
    .ADR3(_n0025),
    .O(\_n0013<28>22/O )
  );
  X_BUF \key2<25>961_G/LUT4_L_BUF  (
    .I(\key2<25>961_G/O ),
    .O(N5635)
  );
  defparam \key2<25>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<25>961_G  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out88 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .O(\key2<25>961_G/O )
  );
  X_BUF \_n0013<26>22/LUT4_L_BUF  (
    .I(\_n0013<26>22/O ),
    .O(_n0013[26])
  );
  defparam \_n0013<26>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<26>22  (
    .ADR0(CHOICE840),
    .ADR1(N5478),
    .ADR2(cipherout2[27]),
    .ADR3(_n0025),
    .O(\_n0013<26>22/O )
  );
  X_BUF \_n0013<24>22/LUT4_L_BUF  (
    .I(\_n0013<24>22/O ),
    .O(_n0013[24])
  );
  defparam \_n0013<24>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<24>22  (
    .ADR0(CHOICE1002),
    .ADR1(N5480),
    .ADR2(N5913),
    .ADR3(_n0025),
    .O(\_n0013<24>22/O )
  );
  X_BUF \key2<37>961_G/LUT4_L_BUF  (
    .I(\key2<37>961_G/O ),
    .O(N5637)
  );
  defparam \key2<37>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<37>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out21 ),
    .O(\key2<37>961_G/O )
  );
  X_BUF \_n0013<22>22/LUT4_L_BUF  (
    .I(\_n0013<22>22/O ),
    .O(_n0013[22])
  );
  defparam \_n0013<22>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<22>22  (
    .ADR0(CHOICE1020),
    .ADR1(N5482),
    .ADR2(cipherout2[23]),
    .ADR3(_n0025),
    .O(\_n0013<22>22/O )
  );
  X_BUF \_n0013<20>22/LUT4_L_BUF  (
    .I(\_n0013<20>22/O ),
    .O(_n0013[20])
  );
  defparam \_n0013<20>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<20>22  (
    .ADR0(CHOICE1011),
    .ADR1(N5484),
    .ADR2(cipherout2[21]),
    .ADR3(_n0025),
    .O(\_n0013<20>22/O )
  );
  X_BUF \_n0013<17>20/LUT4_L_BUF  (
    .I(\_n0013<17>20/O ),
    .O(_n0013[17])
  );
  defparam \_n0013<17>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<17>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1047),
    .ADR2(cipherout2[27]),
    .ADR3(N5017),
    .O(\_n0013<17>20/O )
  );
  X_BUF \_n0013<18>17/LUT4_L_BUF  (
    .I(\_n0013<18>17/O ),
    .O(_n0013[18])
  );
  defparam \_n0013<18>17 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<18>17  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(N5495),
    .ADR3(cipherout2[19]),
    .O(\_n0013<18>17/O )
  );
  X_BUF \_n0013<13>20_SW1/LUT4_L_BUF  (
    .I(\_n0013<13>20_SW1/O ),
    .O(N5432)
  );
  defparam \_n0013<13>20_SW1 .INIT = 16'hECA0;
  X_LUT4 \_n0013<13>20_SW1  (
    .ADR0(data1[14]),
    .ADR1(\state_FFd3-In ),
    .ADR2(N01),
    .ADR3(cipherout2[10]),
    .O(\_n0013<13>20_SW1/O )
  );
  X_BUF \_n0013<16>22/LUT4_L_BUF  (
    .I(\_n0013<16>22/O ),
    .O(_n0013[16])
  );
  defparam \_n0013<16>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<16>22  (
    .ADR0(CHOICE873),
    .ADR1(N5486),
    .ADR2(cipherout2[17]),
    .ADR3(_n0025),
    .O(\_n0013<16>22/O )
  );
  X_BUF \key2<38>961_G/LUT4_L_BUF  (
    .I(\key2<38>961_G/O ),
    .O(N5639)
  );
  defparam \key2<38>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<38>961_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out78 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out40 ),
    .O(\key2<38>961_G/O )
  );
  X_BUF \_n0013<14>22/LUT4_L_BUF  (
    .I(\_n0013<14>22/O ),
    .O(_n0013[14])
  );
  defparam \_n0013<14>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<14>22  (
    .ADR0(CHOICE1038),
    .ADR1(N5448),
    .ADR2(cipherout2[15]),
    .ADR3(_n0025),
    .O(\_n0013<14>22/O )
  );
  X_BUF \_n0013<12>22/LUT4_L_BUF  (
    .I(\_n0013<12>22/O ),
    .O(_n0013[12])
  );
  defparam \_n0013<12>22 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<12>22  (
    .ADR0(CHOICE1029),
    .ADR1(N5488),
    .ADR2(cipherout2[13]),
    .ADR3(_n0025),
    .O(\_n0013<12>22/O )
  );
  X_BUF \key2<3>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<3>133_SW01_G/O ),
    .O(N5641)
  );
  defparam \key2<3>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<3>133_SW01_G  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out74 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out61 ),
    .O(\key2<3>133_SW01_G/O )
  );
  X_BUF \state_FFd3-In1/LUT4_D_BUF  (
    .I(\state_FFd3-In ),
    .O(N5899)
  );
  defparam \state_FFd3-In1 .INIT = 16'hECA0;
  X_LUT4 \state_FFd3-In1  (
    .ADR0(state_FFd4),
    .ADR1(state_FFd2),
    .ADR2(_n0000),
    .ADR3(N5902),
    .O(\state_FFd3-In )
  );
  X_BUF \_n0013<14>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<14>22_SW0/O ),
    .O(N5448)
  );
  defparam \_n0013<14>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<14>22_SW0  (
    .ADR0(data1[2]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[15]),
    .ADR3(N01),
    .O(\_n0013<14>22_SW0/O )
  );
  X_BUF \key2<25>110_SW0/LUT3_L_BUF  (
    .I(\key2<25>110_SW0/O ),
    .O(N5117)
  );
  defparam \key2<25>110_SW0 .INIT = 8'h07;
  X_LUT3 \key2<25>110_SW0  (
    .ADR0(roundsel_2_10),
    .ADR1(N5173),
    .ADR2(CHOICE1134),
    .O(\key2<25>110_SW0/O )
  );
  X_BUF \key2<25>12_SW0_G/LUT3_L_BUF  (
    .I(\key2<25>12_SW0_G/O ),
    .O(N5643)
  );
  defparam \key2<25>12_SW0_G .INIT = 8'hE4;
  X_LUT3 \key2<25>12_SW0_G  (
    .ADR0(roundsel_1_17),
    .ADR1(\key1[8] ),
    .ADR2(\key1[16] ),
    .O(\key2<25>12_SW0_G/O )
  );
  X_BUF \key2<21>1191_G/LUT4_L_BUF  (
    .I(\key2<21>1191_G/O ),
    .O(N5645)
  );
  defparam \key2<21>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<21>1191_G  (
    .ADR0(roundsel_2_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .ADR2(roundsel_3_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .O(\key2<21>1191_G/O )
  );
  X_BUF \key2<33>961_G/LUT4_L_BUF  (
    .I(\key2<33>961_G/O ),
    .O(N5647)
  );
  defparam \key2<33>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<33>961_G  (
    .ADR0(roundsel_3_2),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out80 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out94 ),
    .O(\key2<33>961_G/O )
  );
  X_BUF \_n0013<1>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<1>20_SW0/O ),
    .O(N5033)
  );
  defparam \_n0013<1>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<1>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1945),
    .ADR3(cipherout2[2]),
    .O(\_n0013<1>20_SW0/O )
  );
  X_BUF \key2<13>110_SW0/LUT3_L_BUF  (
    .I(\key2<13>110_SW0/O ),
    .O(N5115)
  );
  defparam \key2<13>110_SW0 .INIT = 8'h07;
  X_LUT3 \key2<13>110_SW0  (
    .ADR0(roundsel[2]),
    .ADR1(N5195),
    .ADR2(CHOICE475),
    .O(\key2<13>110_SW0/O )
  );
  X_BUF \roundsel<2>_mmx_out271_G/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out271_G/O ),
    .O(N5649)
  );
  defparam \roundsel<2>_mmx_out271_G .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out271_G  (
    .ADR0(roundsel_12),
    .ADR1(\key1[50] ),
    .ADR2(\key1[3] ),
    .O(\roundsel<2>_mmx_out271_G/O )
  );
  X_BUF \key2<21>133_SW0/LUT4_L_BUF  (
    .I(\key2<21>133_SW0/O ),
    .O(N5099)
  );
  defparam \key2<21>133_SW0 .INIT = 16'h005D;
  X_LUT4 \key2<21>133_SW0  (
    .ADR0(roundsel_4_5),
    .ADR1(N5131),
    .ADR2(CHOICE970),
    .ADR3(CHOICE980),
    .O(\key2<21>133_SW0/O )
  );
  X_BUF \key2<27>156_SW0/LUT4_L_BUF  (
    .I(\key2<27>156_SW0/O ),
    .O(N5101)
  );
  defparam \key2<27>156_SW0 .INIT = 16'h0705;
  X_LUT4 \key2<27>156_SW0  (
    .ADR0(roundsel_2_12),
    .ADR1(CHOICE1310),
    .ADR2(CHOICE1320),
    .ADR3(N5133),
    .O(\key2<27>156_SW0/O )
  );
  X_BUF \key2<37>110_SW0/LUT3_L_BUF  (
    .I(\key2<37>110_SW0/O ),
    .O(N5119)
  );
  defparam \key2<37>110_SW0 .INIT = 8'h07;
  X_LUT3 \key2<37>110_SW0  (
    .ADR0(roundsel[2]),
    .ADR1(N5175),
    .ADR2(CHOICE1162),
    .O(\key2<37>110_SW0/O )
  );
  X_BUF \key2<28>133_SW0/LUT4_L_BUF  (
    .I(\key2<28>133_SW0/O ),
    .O(N5103)
  );
  defparam \key2<28>133_SW0 .INIT = 16'h0705;
  X_LUT4 \key2<28>133_SW0  (
    .ADR0(roundsel_4_5),
    .ADR1(CHOICE1823),
    .ADR2(CHOICE1833),
    .ADR3(N5135),
    .O(\key2<28>133_SW0/O )
  );
  X_BUF \key2<22>961_G/LUT4_L_BUF  (
    .I(\key2<22>961_G/O ),
    .O(N5651)
  );
  defparam \key2<22>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<22>961_G  (
    .ADR0(roundsel_3_14),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out37 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out33 ),
    .O(\key2<22>961_G/O )
  );
  X_BUF \Ker039/LUT4_D_BUF  (
    .I(N01),
    .O(N5900)
  );
  defparam Ker039_251.INIT = 16'hFFF2;
  X_LUT4 Ker039_251 (
    .ADR0(state_FFd2),
    .ADR1(_n0001),
    .ADR2(CHOICE195),
    .ADR3(CHOICE199),
    .O(N01)
  );
  X_BUF \key2<45>133_SW0/LUT4_L_BUF  (
    .I(\key2<45>133_SW0/O ),
    .O(N5111)
  );
  defparam \key2<45>133_SW0 .INIT = 16'h0705;
  X_LUT4 \key2<45>133_SW0  (
    .ADR0(roundsel_4_9),
    .ADR1(CHOICE1855),
    .ADR2(CHOICE1865),
    .ADR3(N5137),
    .O(\key2<45>133_SW0/O )
  );
  X_BUF \_n0013<29>20_SW0_SW0/LUT4_L_BUF  (
    .I(\_n0013<29>20_SW0_SW0/O ),
    .O(N5151)
  );
  defparam \_n0013<29>20_SW0_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<29>20_SW0_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1954),
    .ADR3(cipherout2[30]),
    .O(\_n0013<29>20_SW0_SW0/O )
  );
  X_BUF \key2<43>110_SW0/LUT3_L_BUF  (
    .I(\key2<43>110_SW0/O ),
    .O(N5121)
  );
  defparam \key2<43>110_SW0 .INIT = 8'h07;
  X_LUT3 \key2<43>110_SW0  (
    .ADR0(roundsel[2]),
    .ADR1(N5177),
    .ADR2(CHOICE1190),
    .O(\key2<43>110_SW0/O )
  );
  X_BUF \_n00001/LUT4_D_BUF  (
    .I(_n0000),
    .O(N5901)
  );
  defparam _n00001.INIT = 16'h8000;
  X_LUT4 _n00001 (
    .ADR0(roundsel_2_10),
    .ADR1(roundsel[1]),
    .ADR2(roundsel_4_5),
    .ADR3(roundsel_3_16),
    .O(_n0000)
  );
  X_BUF \key2<32>12_G/LUT4_L_BUF  (
    .I(\key2<32>12_G/O ),
    .O(N5653)
  );
  defparam \key2<32>12_G .INIT = 16'hA280;
  X_LUT4 \key2<32>12_G  (
    .ADR0(roundsel_2_4),
    .ADR1(roundsel_1_7),
    .ADR2(\key1[13] ),
    .ADR3(\key1[5] ),
    .O(\key2<32>12_G/O )
  );
  X_BUF \_n00011/LUT4_D_BUF  (
    .I(_n0001),
    .O(N5902)
  );
  defparam _n00011.INIT = 16'h0001;
  X_LUT4 _n00011 (
    .ADR0(roundsel[1]),
    .ADR1(roundsel[2]),
    .ADR2(roundsel[4]),
    .ADR3(roundsel[3]),
    .O(_n0001)
  );
  X_BUF \roundsel<1>_mmx_out521/LUT3_D_BUF  (
    .I(\MUX_BLOCK_roundsel<1>_mmx_out52 ),
    .O(N5903)
  );
  defparam \roundsel<1>_mmx_out521 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out521  (
    .ADR0(\key1[59] ),
    .ADR1(\key1[43] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out52 )
  );
  X_BUF \roundsel<1>_mmx_out571/LUT3_D_BUF  (
    .I(\MUX_BLOCK_roundsel<1>_mmx_out57 ),
    .O(N5904)
  );
  defparam \roundsel<1>_mmx_out571 .INIT = 8'hAC;
  X_LUT3 \roundsel<1>_mmx_out571  (
    .ADR0(\key1[26] ),
    .ADR1(\key1[18] ),
    .ADR2(roundsel_1_14),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out57 )
  );
  X_BUF \roundsel<1>_mmx_out621/LUT3_L_BUF  (
    .I(\roundsel<1>_mmx_out621/O ),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out62 )
  );
  defparam \roundsel<1>_mmx_out621 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out621  (
    .ADR0(\key1[60] ),
    .ADR1(\key1[37] ),
    .ADR2(roundsel_1_15),
    .O(\roundsel<1>_mmx_out621/O )
  );
  X_BUF \roundsel<1>_mmx_out631/LUT3_D_BUF  (
    .I(\MUX_BLOCK_roundsel<1>_mmx_out63 ),
    .O(N5905)
  );
  defparam \roundsel<1>_mmx_out631 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out631  (
    .ADR0(\key1[44] ),
    .ADR1(\key1[52] ),
    .ADR2(roundsel_1_9),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out63 )
  );
  X_BUF \roundsel<1>_mmx_out751/LUT3_L_BUF  (
    .I(\roundsel<1>_mmx_out751/O ),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out75 )
  );
  defparam \roundsel<1>_mmx_out751 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out751  (
    .ADR0(\key1[34] ),
    .ADR1(\key1[42] ),
    .ADR2(roundsel_1_5),
    .O(\roundsel<1>_mmx_out751/O )
  );
  X_BUF \roundsel<1>_mmx_out84/LUT3_D_BUF  (
    .I(\MUX_BLOCK_roundsel<1>_mmx_out8 ),
    .O(N5906)
  );
  defparam \roundsel<1>_mmx_out84 .INIT = 8'hCA;
  X_LUT3 \roundsel<1>_mmx_out84  (
    .ADR0(\key1[21] ),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_1_7),
    .O(\MUX_BLOCK_roundsel<1>_mmx_out8 )
  );
  X_BUF \roundsel<2>_mmx_out71_G/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out71_G/O ),
    .O(N5655)
  );
  defparam \roundsel<2>_mmx_out71_G .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out71_G  (
    .ADR0(roundsel_1_16),
    .ADR1(\key1[5] ),
    .ADR2(\key1[21] ),
    .O(\roundsel<2>_mmx_out71_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<7>1/LUT4_D_BUF  (
    .I(cipherout2[8]),
    .O(N5907)
  );
  defparam \c1/Mxor_OUTR_Result<7>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<7>1  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[40]),
    .ADR2(\c1/u4/Mrom_dout_N6 ),
    .ADR3(\c1/u4/Mrom_dout_N7 ),
    .O(cipherout2[8])
  );
  X_BUF \key2<29>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<29>133_SW01_G/O ),
    .O(N5657)
  );
  defparam \key2<29>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<29>133_SW01_G  (
    .ADR0(roundsel_4_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out2 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out85 ),
    .O(\key2<29>133_SW01_G/O )
  );
  X_BUF \key2<41>961_G/LUT4_L_BUF  (
    .I(\key2<41>961_G/O ),
    .O(N5659)
  );
  defparam \key2<41>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<41>961_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out79 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out81 ),
    .O(\key2<41>961_G/O )
  );
  X_BUF \key2<19>761_G/LUT4_L_BUF  (
    .I(\key2<19>761_G/O ),
    .O(N5661)
  );
  defparam \key2<19>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<19>761_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out49 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out32 ),
    .O(\key2<19>761_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<13>1/LUT4_D_BUF  (
    .I(cipherout2[14]),
    .O(N5908)
  );
  defparam \c1/Mxor_OUTR_Result<13>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<13>1  (
    .ADR0(\c1/X[36] ),
    .ADR1(data1[46]),
    .ADR2(\c1/u5/Mrom_dout_N9 ),
    .ADR3(\c1/u5/Mrom_dout_N10 ),
    .O(cipherout2[14])
  );
  X_BUF \c1/Mxor_OUTR_Result<14>1/LUT4_D_BUF  (
    .I(cipherout2[15]),
    .O(N5909)
  );
  defparam \c1/Mxor_OUTR_Result<14>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<14>1  (
    .ADR0(\c1/X[12] ),
    .ADR1(data1[47]),
    .ADR2(\c1/u1/Mrom_dout_N9 ),
    .ADR3(\c1/u1/Mrom_dout_N10 ),
    .O(cipherout2[15])
  );
  X_BUF \roundsel<2>_mmx_out111_G/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out111_G/O ),
    .O(N5663)
  );
  defparam \roundsel<2>_mmx_out111_G .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out111_G  (
    .ADR0(roundsel_1_20),
    .ADR1(\key1[15] ),
    .ADR2(\key1[31] ),
    .O(\roundsel<2>_mmx_out111_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<4>1/LUT4_D_BUF  (
    .I(cipherout2[5]),
    .O(N5910)
  );
  defparam \c1/Mxor_OUTR_Result<4>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<4>1  (
    .ADR0(\c1/X[12] ),
    .ADR1(data1[37]),
    .ADR2(\c1/u1/Mrom_dout_N3 ),
    .ADR3(\c1/u1/Mrom_dout_N4 ),
    .O(cipherout2[5])
  );
  X_BUF \c1/Mxor_OUTR_Result<20>1/LUT4_D_BUF  (
    .I(cipherout2[21]),
    .O(N5911)
  );
  defparam \c1/Mxor_OUTR_Result<20>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<20>1  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[53]),
    .ADR2(\c1/u6/Mrom_dout_N3 ),
    .ADR3(\c1/u6/Mrom_dout_N4 ),
    .O(cipherout2[21])
  );
  X_BUF \c1/Mxor_OUTR_Result<21>1/LUT4_D_BUF  (
    .I(cipherout2[22]),
    .O(N5912)
  );
  defparam \c1/Mxor_OUTR_Result<21>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<21>1  (
    .ADR0(\c1/X[36] ),
    .ADR1(data1[54]),
    .ADR2(\c1/u5/Mrom_dout_N6 ),
    .ADR3(\c1/u5/Mrom_dout_N7 ),
    .O(cipherout2[22])
  );
  X_BUF \c1/Mxor_OUTR_Result<24>1/LUT4_D_BUF  (
    .I(cipherout2[25]),
    .O(N5913)
  );
  defparam \c1/Mxor_OUTR_Result<24>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<24>1  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[57]),
    .ADR2(\c1/u4/Mrom_dout_N0 ),
    .ADR3(\c1/u4/Mrom_dout_N1 ),
    .O(cipherout2[25])
  );
  X_BUF \key2<39>761_G/LUT4_L_BUF  (
    .I(\key2<39>761_G/O ),
    .O(N5665)
  );
  defparam \key2<39>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<39>761_G  (
    .ADR0(roundsel_3_14),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out10 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .O(\key2<39>761_G/O )
  );
  X_BUF \_n0013<11>20/LUT4_L_BUF  (
    .I(\_n0013<11>20/O ),
    .O(_n0013[11])
  );
  defparam \_n0013<11>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<11>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1937),
    .ADR2(cipherout2[18]),
    .ADR3(N5047),
    .O(\_n0013<11>20/O )
  );
  X_BUF \_n0013<31>20_SW0_SW0/LUT4_L_BUF  (
    .I(\_n0013<31>20_SW0_SW0/O ),
    .O(N5193)
  );
  defparam \_n0013<31>20_SW0_SW0 .INIT = 16'hFEEE;
  X_LUT4 \_n0013<31>20_SW0_SW0  (
    .ADR0(CHOICE1964),
    .ADR1(CHOICE1963),
    .ADR2(cipherout2[4]),
    .ADR3(\state_FFd3-In ),
    .O(\_n0013<31>20_SW0_SW0/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<28>1/LUT4_D_BUF  (
    .I(cipherout2[29]),
    .O(N5914)
  );
  defparam \c1/Mxor_OUTR_Result<28>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<28>1  (
    .ADR0(\c1/X[36] ),
    .ADR1(data1[61]),
    .ADR2(\c1/u5/Mrom_dout_N0 ),
    .ADR3(\c1/u5/Mrom_dout_N1 ),
    .O(cipherout2[29])
  );
  X_BUF \c1/Mxor_OUTR_Result<30>1/LUT4_D_BUF  (
    .I(cipherout2[31]),
    .O(N5915)
  );
  defparam \c1/Mxor_OUTR_Result<30>1 .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<30>1  (
    .ADR0(\c1/X[12] ),
    .ADR1(data1[63]),
    .ADR2(\c1/u1/Mrom_dout_N6 ),
    .ADR3(\c1/u1/Mrom_dout_N7 ),
    .O(cipherout2[31])
  );
  X_BUF \c1/Mxor_X_Result<8>1/LUT4_D_BUF  (
    .I(\c1/X[9] ),
    .O(N5916)
  );
  defparam \c1/Mxor_X_Result<8>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<8>1  (
    .ADR0(data1[27]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1437),
    .ADR3(N5093),
    .O(\c1/X[9] )
  );
  X_BUF \c1/Mxor_X_Result<9>1/LUT4_D_BUF  (
    .I(\c1/X[10] ),
    .O(N5917)
  );
  defparam \c1/Mxor_X_Result<9>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<9>1  (
    .ADR0(data1[26]),
    .ADR1(roundsel[4]),
    .ADR2(N5059),
    .ADR3(CHOICE1262),
    .O(\c1/X[10] )
  );
  X_BUF \c1/Mxor_X_Result<10>1/LUT4_D_BUF  (
    .I(\c1/X[11] ),
    .O(N5918)
  );
  defparam \c1/Mxor_X_Result<10>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<10>1  (
    .ADR0(data1[25]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1521),
    .ADR3(N5061),
    .O(\c1/X[11] )
  );
  X_BUF \c1/Mxor_X_Result<13>1/LUT4_D_BUF  (
    .I(\c1/X[14] ),
    .O(N5919)
  );
  defparam \c1/Mxor_X_Result<13>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<13>1  (
    .ADR0(data1[24]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE579),
    .ADR3(N5063),
    .O(\c1/X[14] )
  );
  X_BUF \c1/Mxor_X_Result<14>1/LUT4_D_BUF  (
    .I(\c1/X[15] ),
    .O(N5920)
  );
  defparam \c1/Mxor_X_Result<14>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<14>1  (
    .ADR0(data1[23]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE611),
    .ADR3(N5095),
    .O(\c1/X[15] )
  );
  X_BUF \c1/Mxor_X_Result<16>1/LUT4_D_BUF  (
    .I(\c1/X[17] ),
    .O(N5921)
  );
  defparam \c1/Mxor_X_Result<16>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<16>1  (
    .ADR0(data1[21]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE547),
    .ADR3(N5097),
    .O(\c1/X[17] )
  );
  X_BUF \c1/Mxor_X_Result<19>1/LUT4_D_BUF  (
    .I(\c1/X[20] ),
    .O(N5922)
  );
  defparam \c1/Mxor_X_Result<19>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<19>1  (
    .ADR0(data1[20]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE964),
    .ADR3(N5065),
    .O(\c1/X[20] )
  );
  X_BUF \c1/Mxor_X_Result<21>1/LUT4_D_BUF  (
    .I(\c1/X[22] ),
    .O(N5923)
  );
  defparam \c1/Mxor_X_Result<21>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<21>1  (
    .ADR0(data1[18]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE936),
    .ADR3(N5067),
    .O(\c1/X[22] )
  );
  X_BUF \c1/Mxor_X_Result<22>1/LUT4_D_BUF  (
    .I(\c1/X[23] ),
    .O(N5924)
  );
  defparam \c1/Mxor_X_Result<22>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<22>1  (
    .ADR0(data1[17]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE908),
    .ADR3(N5069),
    .O(\c1/X[23] )
  );
  X_BUF \c1/Mxor_X_Result<28>1/LUT4_D_BUF  (
    .I(\c1/X[29] ),
    .O(N5925)
  );
  defparam \c1/Mxor_X_Result<28>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<28>1  (
    .ADR0(data1[13]),
    .ADR1(roundsel[3]),
    .ADR2(CHOICE1553),
    .ADR3(N5071),
    .O(\c1/X[29] )
  );
  X_BUF \c1/Mxor_X_Result<32>1/LUT4_D_BUF  (
    .I(\c1/X[33] ),
    .O(N5926)
  );
  defparam \c1/Mxor_X_Result<32>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<32>1  (
    .ADR0(data1[11]),
    .ADR1(roundsel_4_5),
    .ADR2(CHOICE1493),
    .ADR3(N5073),
    .O(\c1/X[33] )
  );
  X_BUF \c1/Mxor_X_Result<33>1/LUT4_D_BUF  (
    .I(\c1/X[34] ),
    .O(N5927)
  );
  defparam \c1/Mxor_X_Result<33>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<33>1  (
    .ADR0(data1[10]),
    .ADR1(roundsel_4_5),
    .ADR2(N5075),
    .ADR3(CHOICE1234),
    .O(\c1/X[34] )
  );
  X_BUF \c1/Mxor_X_Result<34>1/LUT4_D_BUF  (
    .I(\c1/X[35] ),
    .O(N5928)
  );
  defparam \c1/Mxor_X_Result<34>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<34>1  (
    .ADR0(data1[9]),
    .ADR1(roundsel_4_5),
    .ADR2(CHOICE1304),
    .ADR3(N5105),
    .O(\c1/X[35] )
  );
  X_BUF \c1/Mxor_X_Result<37>1/LUT4_D_BUF  (
    .I(\c1/X[38] ),
    .O(N5929)
  );
  defparam \c1/Mxor_X_Result<37>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<37>1  (
    .ADR0(data1[8]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1817),
    .ADR3(N5077),
    .O(\c1/X[38] )
  );
  X_BUF \c1/Mxor_X_Result<38>1/LUT4_D_BUF  (
    .I(\c1/X[39] ),
    .O(N5930)
  );
  defparam \c1/Mxor_X_Result<38>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<38>1  (
    .ADR0(data1[7]),
    .ADR1(roundsel[4]),
    .ADR2(N5107),
    .ADR3(CHOICE1609),
    .O(\c1/X[39] )
  );
  X_BUF \c1/Mxor_X_Result<39>1/LUT4_D_BUF  (
    .I(\c1/X[40] ),
    .O(N5931)
  );
  defparam \c1/Mxor_X_Result<39>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<39>1  (
    .ADR0(data1[6]),
    .ADR1(roundsel[3]),
    .ADR2(CHOICE1705),
    .ADR3(N5109),
    .O(\c1/X[40] )
  );
  X_BUF \c1/Mxor_X_Result<40>1/LUT4_D_BUF  (
    .I(\c1/X[41] ),
    .O(N5932)
  );
  defparam \c1/Mxor_X_Result<40>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<40>1  (
    .ADR0(data1[5]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1465),
    .ADR3(N5079),
    .O(\c1/X[41] )
  );
  X_BUF \c1/Mxor_X_Result<43>1/LUT4_D_BUF  (
    .I(\c1/X[44] ),
    .O(N5933)
  );
  defparam \c1/Mxor_X_Result<43>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<43>1  (
    .ADR0(data1[4]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1789),
    .ADR3(N5081),
    .O(\c1/X[44] )
  );
  X_BUF \c1/Mxor_X_Result<45>1/LUT4_D_BUF  (
    .I(\c1/X[46] ),
    .O(N5934)
  );
  defparam \c1/Mxor_X_Result<45>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<45>1  (
    .ADR0(data1[2]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1913),
    .ADR3(N5113),
    .O(\c1/X[46] )
  );
  X_BUF \c1/Mxor_X_Result<46>1/LUT4_D_BUF  (
    .I(\c1/X[47] ),
    .O(N5935)
  );
  defparam \c1/Mxor_X_Result<46>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<46>1  (
    .ADR0(data1[1]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1377),
    .ADR3(N5083),
    .O(\c1/X[47] )
  );
  X_BUF \c1/Mxor_X_Result<2>1/LUT4_D_BUF  (
    .I(\c1/X[3] ),
    .O(N5936)
  );
  defparam \c1/Mxor_X_Result<2>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<2>1  (
    .ADR0(data1[31]),
    .ADR1(roundsel[2]),
    .ADR2(N5085),
    .ADR3(CHOICE1585),
    .O(\c1/X[3] )
  );
  X_BUF \c1/Mxor_X_Result<1>1/LUT4_D_BUF  (
    .I(\c1/X[2] ),
    .O(N5937)
  );
  defparam \c1/Mxor_X_Result<1>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<1>1  (
    .ADR0(data1[32]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1733),
    .ADR3(N5087),
    .O(\c1/X[2] )
  );
  X_BUF \c1/Mxor_X_Result<3>1/LUT4_D_BUF  (
    .I(\c1/X[4] ),
    .O(N5938)
  );
  defparam \c1/Mxor_X_Result<3>1 .INIT = 16'h55A6;
  X_LUT4 \c1/Mxor_X_Result<3>1  (
    .ADR0(data1[30]),
    .ADR1(roundsel[4]),
    .ADR2(N5089),
    .ADR3(CHOICE1761),
    .O(\c1/X[4] )
  );
  X_BUF \key2<31>761_G/LUT4_L_BUF  (
    .I(\key2<31>761_G/O ),
    .O(N5667)
  );
  defparam \key2<31>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<31>761_G  (
    .ADR0(roundsel_3_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out81 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out95 ),
    .O(\key2<31>761_G/O )
  );
  X_BUF \c1/Mxor_X_Result<4>1/LUT4_D_BUF  (
    .I(\c1/X[5] ),
    .O(N5939)
  );
  defparam \c1/Mxor_X_Result<4>1 .INIT = 16'h5A56;
  X_LUT4 \c1/Mxor_X_Result<4>1  (
    .ADR0(data1[29]),
    .ADR1(roundsel[4]),
    .ADR2(CHOICE1405),
    .ADR3(N5091),
    .O(\c1/X[5] )
  );
  X_BUF \key2<4>961_G/LUT4_L_BUF  (
    .I(\key2<4>961_G/O ),
    .O(N5669)
  );
  defparam \key2<4>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<4>961_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out41 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out50 ),
    .O(\key2<4>961_G/O )
  );
  X_BUF \_n0013<23>20/LUT4_L_BUF  (
    .I(\_n0013<23>20/O ),
    .O(_n0013[23])
  );
  defparam \_n0013<23>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<23>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1277),
    .ADR2(cipherout2[3]),
    .ADR3(N5035),
    .O(\_n0013<23>20/O )
  );
  X_BUF \key2<47>961_G/LUT4_L_BUF  (
    .I(\key2<47>961_G/O ),
    .O(N5671)
  );
  defparam \key2<47>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<47>961_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out77 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out31 ),
    .O(\key2<47>961_G/O )
  );
  X_BUF \key2<17>25_SW0/LUT4_L_BUF  (
    .I(\key2<17>25_SW0/O ),
    .O(N5141)
  );
  defparam \key2<17>25_SW0 .INIT = 16'hFF53;
  X_LUT4 \key2<17>25_SW0  (
    .ADR0(\key1[3] ),
    .ADR1(\key1[50] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_23),
    .O(\key2<17>25_SW0/O )
  );
  X_BUF \key2<44>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<44>110_SW01_G/O ),
    .O(N5673)
  );
  defparam \key2<44>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<44>110_SW01_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out1 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out95 ),
    .O(\key2<44>110_SW01_G/O )
  );
  X_BUF \key2<34>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<34>110_SW01_G/O ),
    .O(N5675)
  );
  defparam \key2<34>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<34>110_SW01_G  (
    .ADR0(roundsel_3_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out18 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out20 ),
    .O(\key2<34>110_SW01_G/O )
  );
  X_BUF \key2<43>961_G/LUT4_L_BUF  (
    .I(\key2<43>961_G/O ),
    .O(N5677)
  );
  defparam \key2<43>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<43>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out55 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out3 ),
    .O(\key2<43>961_G/O )
  );
  X_BUF \c1/Mxor_X_Result<7>11_G/LUT3_L_BUF  (
    .I(\c1/Mxor_X_Result<7>11_G/O ),
    .O(N5679)
  );
  defparam \c1/Mxor_X_Result<7>11_G .INIT = 8'h56;
  X_LUT3 \c1/Mxor_X_Result<7>11_G  (
    .ADR0(data1[28]),
    .ADR1(CHOICE1621),
    .ADR2(CHOICE1615),
    .O(\c1/Mxor_X_Result<7>11_G/O )
  );
  X_BUF \key2<35>761_G/LUT4_L_BUF  (
    .I(\key2<35>761_G/O ),
    .O(N5681)
  );
  defparam \key2<35>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<35>761_G  (
    .ADR0(roundsel_3_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out86 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out20 ),
    .O(\key2<35>761_G/O )
  );
  X_BUF \key2<45>471_G/LUT4_L_BUF  (
    .I(\key2<45>471_G/O ),
    .O(N5683)
  );
  defparam \key2<45>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<45>471_G  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[48] ),
    .ADR2(roundsel_4_1),
    .ADR3(\key1[15] ),
    .O(\key2<45>471_G/O )
  );
  X_BUF \_n0013<3>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<3>20_SW0/O ),
    .O(N5434)
  );
  defparam \_n0013<3>20_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<3>20_SW0  (
    .ADR0(data1[4]),
    .ADR1(\state_FFd3-In ),
    .ADR2(N01),
    .ADR3(cipherout2[17]),
    .O(\_n0013<3>20_SW0/O )
  );
  X_BUF \key2<6>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<6>110_SW01_G/O ),
    .O(N5685)
  );
  defparam \key2<6>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<6>110_SW01_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out70 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .O(\key2<6>110_SW01_G/O )
  );
  X_BUF \key2<34>961_G/LUT4_L_BUF  (
    .I(\key2<34>961_G/O ),
    .O(N5687)
  );
  defparam \key2<34>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<34>961_G  (
    .ADR0(roundsel_3_8),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out94 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out ),
    .O(\key2<34>961_G/O )
  );
  X_BUF \key2<6>961_G/LUT4_L_BUF  (
    .I(\key2<6>961_G/O ),
    .O(N5689)
  );
  defparam \key2<6>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<6>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out39 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out73 ),
    .O(\key2<6>961_G/O )
  );
  X_BUF \key2<35>90_SW01_G/LUT3_L_BUF  (
    .I(\key2<35>90_SW01_G/O ),
    .O(N5691)
  );
  defparam \key2<35>90_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<35>90_SW01_G  (
    .ADR0(roundsel_3_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out76 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out10 ),
    .O(\key2<35>90_SW01_G/O )
  );
  X_BUF \key2<30>1181_G/LUT4_L_BUF  (
    .I(\key2<30>1181_G/O ),
    .O(N5693)
  );
  defparam \key2<30>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<30>1181_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out95 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out90 ),
    .O(\key2<30>1181_G/O )
  );
  X_BUF \key2<17>471_G/LUT4_L_BUF  (
    .I(\key2<17>471_G/O ),
    .O(N5695)
  );
  defparam \key2<17>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<17>471_G  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[2] ),
    .ADR2(roundsel_3_1),
    .ADR3(\key1[34] ),
    .O(\key2<17>471_G/O )
  );
  X_BUF \key2<18>961_G/LUT4_L_BUF  (
    .I(\key2<18>961_G/O ),
    .O(N5697)
  );
  defparam \key2<18>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<18>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out50 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out52 ),
    .O(\key2<18>961_G/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_321/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_321/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_32 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_321 .INIT = 16'hE16A;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_321  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_321/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_341/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_341/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_34 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_341 .INIT = 16'h781D;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_341  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_341/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_381/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_381/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_38 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_381 .INIT = 16'hC996;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_381  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[35] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_381/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_mux_f5_18/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_mux_f5_18/O ),
    .O(\c1/u5/Mrom_dout_N3 )
  );
  defparam \c1/u5/Mrom_dout_inst_mux_f5_18 .INIT = 16'hF690;
  X_LUT4 \c1/u5/Mrom_dout_inst_mux_f5_18  (
    .ADR0(data1[13]),
    .ADR1(\key2[31] ),
    .ADR2(\c1/u5/Mrom_dout_inst_lut4_36 ),
    .ADR3(\c1/u5/Mrom_dout_inst_lut4_37 ),
    .O(\c1/u5/Mrom_dout_inst_mux_f5_18/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_401/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_401/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_40 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_401 .INIT = 16'h7A49;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_401  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[35] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_401/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_421/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_421/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_42 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_421 .INIT = 16'hA54E;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_421  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[34] ),
    .ADR3(\c1/X[35] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_421/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_441/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_441/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_44 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_441 .INIT = 16'h994B;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_441  (
    .ADR0(\c1/X[33] ),
    .ADR1(\c1/X[32] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_441/O )
  );
  X_BUF \c1/u5/Mrom_dout_inst_lut4_461/LUT4_L_BUF  (
    .I(\c1/u5/Mrom_dout_inst_lut4_461/O ),
    .O(\c1/u5/Mrom_dout_inst_lut4_46 )
  );
  defparam \c1/u5/Mrom_dout_inst_lut4_461 .INIT = 16'h6687;
  X_LUT4 \c1/u5/Mrom_dout_inst_lut4_461  (
    .ADR0(\c1/X[32] ),
    .ADR1(\c1/X[33] ),
    .ADR2(\c1/X[35] ),
    .ADR3(\c1/X[34] ),
    .O(\c1/u5/Mrom_dout_inst_lut4_461/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<16>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<16>11_G/O ),
    .O(N5699)
  );
  defparam \c1/Mxor_OUTR_Result<16>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<16>11_G  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[49]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_85 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_87 ),
    .O(\c1/Mxor_OUTR_Result<16>11_G/O )
  );
  X_BUF \key2<42>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<42>110_SW01_G/O ),
    .O(N5701)
  );
  defparam \key2<42>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<42>110_SW01_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out92 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out21 ),
    .O(\key2<42>110_SW01_G/O )
  );
  X_BUF \key2<40>90_SW01_G/LUT3_L_BUF  (
    .I(\key2<40>90_SW01_G/O ),
    .O(N5703)
  );
  defparam \key2<40>90_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<40>90_SW01_G  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out11 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out9 ),
    .O(\key2<40>90_SW01_G/O )
  );
  X_BUF \key2<21>471_G/LUT4_L_BUF  (
    .I(\key2<21>471_G/O ),
    .O(N5705)
  );
  defparam \key2<21>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<21>471_G  (
    .ADR0(roundsel_2_4),
    .ADR1(\key1[20] ),
    .ADR2(roundsel_4_2),
    .ADR3(\key1[52] ),
    .O(\key2<21>471_G/O )
  );
  X_BUF \key2<24>1181_G/LUT4_L_BUF  (
    .I(\key2<24>1181_G/O ),
    .O(N5707)
  );
  defparam \key2<24>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<24>1181_G  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out25 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out26 ),
    .O(\key2<24>1181_G/O )
  );
  X_BUF \key2<48>961_G/LUT4_L_BUF  (
    .I(\key2<48>961_G/O ),
    .O(N5709)
  );
  defparam \key2<48>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<48>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out23 ),
    .O(\key2<48>961_G/O )
  );
  X_BUF \key2<36>1181_G/LUT4_L_BUF  (
    .I(\key2<36>1181_G/O ),
    .O(N5711)
  );
  defparam \key2<36>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<36>1181_G  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out20 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out5 ),
    .O(\key2<36>1181_G/O )
  );
  X_BUF \key2<23>1181_G/LUT4_L_BUF  (
    .I(\key2<23>1181_G/O ),
    .O(N5713)
  );
  defparam \key2<23>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<23>1181_G  (
    .ADR0(roundsel_2_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out28 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out29 ),
    .O(\key2<23>1181_G/O )
  );
  X_BUF \key2<48>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<48>110_SW01_G/O ),
    .O(N5715)
  );
  defparam \key2<48>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<48>110_SW01_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out64 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out40 ),
    .O(\key2<48>110_SW01_G/O )
  );
  X_BUF \c1/Mxor_X_Result<0>11_G/LUT3_L_BUF  (
    .I(\c1/Mxor_X_Result<0>11_G/O ),
    .O(N5717)
  );
  defparam \c1/Mxor_X_Result<0>11_G .INIT = 8'h56;
  X_LUT3 \c1/Mxor_X_Result<0>11_G  (
    .ADR0(data1[1]),
    .ADR1(CHOICE1086),
    .ADR2(CHOICE1080),
    .O(\c1/Mxor_X_Result<0>11_G/O )
  );
  X_BUF \key2<1>271_G/LUT4_L_BUF  (
    .I(\key2<1>271_G/O ),
    .O(N5719)
  );
  defparam \key2<1>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<1>271_G  (
    .ADR0(roundsel_3_16),
    .ADR1(\key1[36] ),
    .ADR2(roundsel[2]),
    .ADR3(\key1[2] ),
    .O(\key2<1>271_G/O )
  );
  X_BUF \key2<44>961_G/LUT4_L_BUF  (
    .I(\key2<44>961_G/O ),
    .O(N5721)
  );
  defparam \key2<44>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<44>961_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out40 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out93 ),
    .O(\key2<44>961_G/O )
  );
  X_BUF \key2<18>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<18>110_SW01_G/O ),
    .O(N5723)
  );
  defparam \key2<18>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<18>110_SW01_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out58 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out25 ),
    .O(\key2<18>110_SW01_G/O )
  );
  X_BUF \key2<36>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<36>133_SW01_G/O ),
    .O(N5725)
  );
  defparam \key2<36>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<36>133_SW01_G  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out16 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .O(\key2<36>133_SW01_G/O )
  );
  X_BUF \key2<16>271_G/LUT4_L_BUF  (
    .I(\key2<16>271_G/O ),
    .O(N5727)
  );
  defparam \key2<16>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<16>271_G  (
    .ADR0(roundsel_3_8),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[28] ),
    .O(\key2<16>271_G/O )
  );
  X_BUF \c1/Mxor_X_Result<25>11_G/LUT3_L_BUF  (
    .I(\c1/Mxor_X_Result<25>11_G/O ),
    .O(N5729)
  );
  defparam \c1/Mxor_X_Result<25>11_G .INIT = 8'h56;
  X_LUT3 \c1/Mxor_X_Result<25>11_G  (
    .ADR0(data1[16]),
    .ADR1(CHOICE1645),
    .ADR2(CHOICE1639),
    .O(\c1/Mxor_X_Result<25>11_G/O )
  );
  X_BUF \key2<14>1181_G/LUT4_L_BUF  (
    .I(\key2<14>1181_G/O ),
    .O(N5731)
  );
  defparam \key2<14>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<14>1181_G  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out24 ),
    .O(\key2<14>1181_G/O )
  );
  X_BUF \key2<12>761_G/LUT4_L_BUF  (
    .I(\key2<12>761_G/O ),
    .O(N5733)
  );
  defparam \key2<12>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<12>761_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out61 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .O(\key2<12>761_G/O )
  );
  X_BUF \c1/u3/Mrom_dout_inst_lut4_781/LUT4_L_BUF  (
    .I(\c1/u3/Mrom_dout_inst_lut4_781/O ),
    .O(\c1/u3/Mrom_dout_inst_lut4_78 )
  );
  defparam \c1/u3/Mrom_dout_inst_lut4_781 .INIT = 16'h619B;
  X_LUT4 \c1/u3/Mrom_dout_inst_lut4_781  (
    .ADR0(\c1/X[22] ),
    .ADR1(\c1/X[20] ),
    .ADR2(\c1/X[21] ),
    .ADR3(\c1/X[23] ),
    .O(\c1/u3/Mrom_dout_inst_lut4_781/O )
  );
  X_BUF \key2<8>61_G/LUT3_L_BUF  (
    .I(\key2<8>61_G/O ),
    .O(N5735)
  );
  defparam \key2<8>61_G .INIT = 8'hE4;
  X_LUT3 \key2<8>61_G  (
    .ADR0(roundsel_12),
    .ADR1(\key1[11] ),
    .ADR2(\key1[27] ),
    .O(\key2<8>61_G/O )
  );
  X_BUF \c1/u3/Mrom_dout_inst_mux_f5_38/LUT4_L_BUF  (
    .I(\c1/u3/Mrom_dout_inst_mux_f5_38/O ),
    .O(\c1/u3/Mrom_dout_N9 )
  );
  defparam \c1/u3/Mrom_dout_inst_mux_f5_38 .INIT = 16'hF690;
  X_LUT4 \c1/u3/Mrom_dout_inst_mux_f5_38  (
    .ADR0(data1[21]),
    .ADR1(\key2[19] ),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_76 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_72 ),
    .O(\c1/u3/Mrom_dout_inst_mux_f5_38/O )
  );
  X_BUF \key2<13>961_G/LUT4_L_BUF  (
    .I(\key2<13>961_G/O ),
    .O(N5737)
  );
  defparam \key2<13>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<13>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out28 ),
    .O(\key2<13>961_G/O )
  );
  X_BUF \key2<19>90_SW0/LUT2_L_BUF  (
    .I(\key2<19>90_SW0/O ),
    .O(N5181)
  );
  defparam \key2<19>90_SW0 .INIT = 4'h1;
  X_LUT2 \key2<19>90_SW0  (
    .ADR0(CHOICE851),
    .ADR1(CHOICE849),
    .O(\key2<19>90_SW0/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<2>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<2>11_G/O ),
    .O(N5739)
  );
  defparam \c1/Mxor_OUTR_Result<2>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<2>11_G  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[35]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_89 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_91 ),
    .O(\c1/Mxor_OUTR_Result<2>11_G/O )
  );
  X_BUF \key2<9>471_G/LUT4_L_BUF  (
    .I(\key2<9>471_G/O ),
    .O(N5741)
  );
  defparam \key2<9>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<9>471_G  (
    .ADR0(roundsel_3_7),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[37] ),
    .O(\key2<9>471_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<1>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<1>11_G/O ),
    .O(N5743)
  );
  defparam \c1/Mxor_OUTR_Result<1>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<1>11_G  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[34]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_109 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_111 ),
    .O(\c1/Mxor_OUTR_Result<1>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<9>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<9>11_G/O ),
    .O(N5745)
  );
  defparam \c1/Mxor_OUTR_Result<9>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<9>11_G  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[42]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_105 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_107 ),
    .O(\c1/Mxor_OUTR_Result<9>11_G/O )
  );
  X_BUF \key2<38>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<38>110_SW01_G/O ),
    .O(N5747)
  );
  defparam \key2<38>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<38>110_SW01_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out17 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out81 ),
    .O(\key2<38>110_SW01_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<15>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<15>11_G/O ),
    .O(N5749)
  );
  defparam \c1/Mxor_OUTR_Result<15>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<15>11_G  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[48]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_101 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_103 ),
    .O(\c1/Mxor_OUTR_Result<15>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<8>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<8>11_G/O ),
    .O(N5751)
  );
  defparam \c1/Mxor_OUTR_Result<8>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<8>11_G  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[41]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_81 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_83 ),
    .O(\c1/Mxor_OUTR_Result<8>11_G/O )
  );
  X_BUF \key2<41>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<41>110_SW01_G/O ),
    .O(N5753)
  );
  defparam \key2<41>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<41>110_SW01_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out8 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out85 ),
    .O(\key2<41>110_SW01_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<26>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<26>11_G/O ),
    .O(N5755)
  );
  defparam \c1/Mxor_OUTR_Result<26>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<26>11_G  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[59]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_93 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_95 ),
    .O(\c1/Mxor_OUTR_Result<26>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<29>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<29>11_G/O ),
    .O(N5757)
  );
  defparam \c1/Mxor_OUTR_Result<29>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<29>11_G  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[62]),
    .ADR2(\c1/u4/Mrom_dout_inst_lut4_61 ),
    .ADR3(\c1/u4/Mrom_dout_inst_lut4_63 ),
    .O(\c1/Mxor_OUTR_Result<29>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<22>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<22>11_G/O ),
    .O(N5759)
  );
  defparam \c1/Mxor_OUTR_Result<22>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<22>11_G  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[55]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_73 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_75 ),
    .O(\c1/Mxor_OUTR_Result<22>11_G/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_lut4_1141/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_lut4_1141/O ),
    .O(\c1/u1/Mrom_dout_inst_lut4_114 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1141 .INIT = 16'hD1AA;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1141  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_1141/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_mux_f5_56/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_mux_f5_56/O ),
    .O(\c1/u1/Mrom_dout_N0 )
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_56 .INIT = 16'hF690;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_56  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/u1/Mrom_dout_inst_lut4_112 ),
    .ADR3(\c1/u1/Mrom_dout_inst_lut4_113 ),
    .O(\c1/u1/Mrom_dout_inst_mux_f5_56/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_lut4_1161/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_lut4_1161/O ),
    .O(\c1/u1/Mrom_dout_inst_lut4_116 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1161 .INIT = 16'h8679;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1161  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_1161/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_lut4_1181/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_lut4_1181/O ),
    .O(\c1/u1/Mrom_dout_inst_lut4_118 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1181 .INIT = 16'hE81E;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1181  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_1181/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_lut4_1201/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_lut4_1201/O ),
    .O(\c1/u1/Mrom_dout_inst_lut4_120 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1201 .INIT = 16'h3C99;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1201  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_1201/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_lut4_1221/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_lut4_1221/O ),
    .O(\c1/u1/Mrom_dout_inst_lut4_122 )
  );
  defparam \c1/u1/Mrom_dout_inst_lut4_1221 .INIT = 16'h8B66;
  X_LUT4 \c1/u1/Mrom_dout_inst_lut4_1221  (
    .ADR0(\c1/X[9] ),
    .ADR1(\c1/X[8] ),
    .ADR2(\c1/X[10] ),
    .ADR3(\c1/X[11] ),
    .O(\c1/u1/Mrom_dout_inst_lut4_1221/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_mux_f5_62_SW1/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_mux_f5_62_SW1/O ),
    .O(N5187)
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_62_SW1 .INIT = 16'h6609;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_62_SW1  (
    .ADR0(data1[29]),
    .ADR1(\key2[7] ),
    .ADR2(\c1/X[11] ),
    .ADR3(\c1/X[10] ),
    .O(\c1/u1/Mrom_dout_inst_mux_f5_62_SW1/O )
  );
  X_BUF \c1/u1/Mrom_dout_inst_mux_f5_63_SW1/LUT4_L_BUF  (
    .I(\c1/u1/Mrom_dout_inst_mux_f5_63_SW1/O ),
    .O(N5184)
  );
  defparam \c1/u1/Mrom_dout_inst_mux_f5_63_SW1 .INIT = 16'hDE69;
  X_LUT4 \c1/u1/Mrom_dout_inst_mux_f5_63_SW1  (
    .ADR0(data1[29]),
    .ADR1(\c1/X[8] ),
    .ADR2(\key2[7] ),
    .ADR3(\c1/X[10] ),
    .O(\c1/u1/Mrom_dout_inst_mux_f5_63_SW1/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<12>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<12>11_G/O ),
    .O(N5763)
  );
  defparam \c1/Mxor_OUTR_Result<12>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<12>11_G  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[45]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_69 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_71 ),
    .O(\c1/Mxor_OUTR_Result<12>11_G/O )
  );
  X_BUF \key2<12>90_SW0_G/LUT3_L_BUF  (
    .I(\key2<12>90_SW0_G/O ),
    .O(N5765)
  );
  defparam \key2<12>90_SW0_G .INIT = 8'h27;
  X_LUT3 \key2<12>90_SW0_G  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out71 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out32 ),
    .O(\key2<12>90_SW0_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<6>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<6>11_G/O ),
    .O(N5767)
  );
  defparam \c1/Mxor_OUTR_Result<6>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<6>11_G  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[39]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_65 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_67 ),
    .O(\c1/Mxor_OUTR_Result<6>11_G/O )
  );
  X_BUF \key2<46>471_G/LUT4_L_BUF  (
    .I(\key2<46>471_G/O ),
    .O(N5769)
  );
  defparam \key2<46>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<46>471_G  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[64] ),
    .O(\key2<46>471_G/O )
  );
  X_BUF \_n0013<48>21/LUT3_L_BUF  (
    .I(\_n0013<48>21/O ),
    .O(_n0013[48])
  );
  defparam \_n0013<48>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<48>21  (
    .ADR0(CHOICE95),
    .ADR1(data1[49]),
    .ADR2(N01),
    .O(\_n0013<48>21/O )
  );
  X_BUF \_n0013<28>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<28>22_SW0/O ),
    .O(N5446)
  );
  defparam \_n0013<28>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<28>22_SW0  (
    .ADR0(data1[12]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[29]),
    .ADR3(N01),
    .O(\_n0013<28>22_SW0/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<27>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<27>11_G/O ),
    .O(N5771)
  );
  defparam \c1/Mxor_OUTR_Result<27>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<27>11_G  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[60]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_1 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_3 ),
    .O(\c1/Mxor_OUTR_Result<27>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<11>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<11>11_G/O ),
    .O(N5773)
  );
  defparam \c1/Mxor_OUTR_Result<11>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<11>11_G  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[44]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_13 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_15 ),
    .O(\c1/Mxor_OUTR_Result<11>11_G/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<23>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<23>11_G/O ),
    .O(N5775)
  );
  defparam \c1/Mxor_OUTR_Result<23>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<23>11_G  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[56]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_97 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_99 ),
    .O(\c1/Mxor_OUTR_Result<23>11_G/O )
  );
  X_BUF \_n0013<42>5/LUT4_L_BUF  (
    .I(\_n0013<42>5/O ),
    .O(CHOICE19)
  );
  defparam \_n0013<42>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<42>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[22]),
    .ADR2(state_FFd8),
    .ADR3(datain_43_IBUF),
    .O(\_n0013<42>5/O )
  );
  X_BUF \_n0013<47>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<47>22_SW0/O ),
    .O(N5470)
  );
  defparam \_n0013<47>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<47>22_SW0  (
    .ADR0(data1[16]),
    .ADR1(_n0025),
    .ADR2(data1[48]),
    .ADR3(N01),
    .O(\_n0013<47>22_SW0/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<10>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<10>11_G/O ),
    .O(N5777)
  );
  defparam \c1/Mxor_OUTR_Result<10>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<10>11_G  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[43]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_25 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_27 ),
    .O(\c1/Mxor_OUTR_Result<10>11_G/O )
  );
  X_BUF \key2<8>271_G/LUT4_L_BUF  (
    .I(\key2<8>271_G/O ),
    .O(N5779)
  );
  defparam \key2<8>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<8>271_G  (
    .ADR0(roundsel_3_8),
    .ADR1(\key1[52] ),
    .ADR2(roundsel_23),
    .ADR3(\key1[18] ),
    .O(\key2<8>271_G/O )
  );
  X_BUF \_n0013<46>5/LUT4_L_BUF  (
    .I(\_n0013<46>5/O ),
    .O(CHOICE100)
  );
  defparam \_n0013<46>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<46>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[54]),
    .ADR2(state_FFd8),
    .ADR3(datain_47_IBUF),
    .O(\_n0013<46>5/O )
  );
  X_BUF \_n0013<34>14/LUT3_L_BUF  (
    .I(\_n0013<34>14/O ),
    .O(CHOICE158)
  );
  defparam \_n0013<34>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<34>14  (
    .ADR0(CHOICE156),
    .ADR1(data1[21]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<34>14/O )
  );
  X_BUF \_n0013<42>14/LUT3_L_BUF  (
    .I(\_n0013<42>14/O ),
    .O(CHOICE23)
  );
  defparam \_n0013<42>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<42>14  (
    .ADR0(CHOICE21),
    .ADR1(data1[22]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<42>14/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<5>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<5>11_G/O ),
    .O(N5781)
  );
  defparam \c1/Mxor_OUTR_Result<5>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<5>11_G  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[38]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_5 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_7 ),
    .O(\c1/Mxor_OUTR_Result<5>11_G/O )
  );
  X_BUF \_n0013<42>21/LUT3_L_BUF  (
    .I(\_n0013<42>21/O ),
    .O(_n0013[42])
  );
  defparam \_n0013<42>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<42>21  (
    .ADR0(CHOICE23),
    .ADR1(data1[43]),
    .ADR2(N01),
    .O(\_n0013<42>21/O )
  );
  X_BUF \_n0013<34>21/LUT3_L_BUF  (
    .I(\_n0013<34>21/O ),
    .O(_n0013[34])
  );
  defparam \_n0013<34>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<34>21  (
    .ADR0(CHOICE158),
    .ADR1(data1[35]),
    .ADR2(N01),
    .O(\_n0013<34>21/O )
  );
  X_BUF \key2<40>761_G/LUT4_L_BUF  (
    .I(\key2<40>761_G/O ),
    .O(N5783)
  );
  defparam \key2<40>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<40>761_G  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out85 ),
    .ADR2(roundsel_3_13),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out88 ),
    .O(\key2<40>761_G/O )
  );
  X_BUF \_n0013<46>14/LUT3_L_BUF  (
    .I(\_n0013<46>14/O ),
    .O(CHOICE104)
  );
  defparam \_n0013<46>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<46>14  (
    .ADR0(CHOICE102),
    .ADR1(data1[6]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<46>14/O )
  );
  X_BUF \_n0013<30>1/LUT2_L_BUF  (
    .I(\_n0013<30>1/O ),
    .O(CHOICE819)
  );
  defparam \_n0013<30>1 .INIT = 4'h8;
  X_LUT2 \_n0013<30>1  (
    .ADR0(data1[31]),
    .ADR1(N01),
    .O(\_n0013<30>1/O )
  );
  X_BUF \_n0013<62>5/LUT4_L_BUF  (
    .I(\_n0013<62>5/O ),
    .O(CHOICE28)
  );
  defparam \_n0013<62>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<62>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[50]),
    .ADR2(state_FFd8),
    .ADR3(datain_63_IBUF),
    .O(\_n0013<62>5/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<18>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<18>11_G/O ),
    .O(N5785)
  );
  defparam \c1/Mxor_OUTR_Result<18>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<18>11_G  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[51]),
    .ADR2(\c1/u4/Mrom_dout_inst_lut4_53 ),
    .ADR3(\c1/u4/Mrom_dout_inst_lut4_55 ),
    .O(\c1/Mxor_OUTR_Result<18>11_G/O )
  );
  X_BUF \_n0013<46>21/LUT3_L_BUF  (
    .I(\_n0013<46>21/O ),
    .O(_n0013[46])
  );
  defparam \_n0013<46>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<46>21  (
    .ADR0(CHOICE104),
    .ADR1(data1[47]),
    .ADR2(N01),
    .O(\_n0013<46>21/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<0>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<0>11_G/O ),
    .O(N5787)
  );
  defparam \c1/Mxor_OUTR_Result<0>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<0>11_G  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[33]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_17 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_19 ),
    .O(\c1/Mxor_OUTR_Result<0>11_G/O )
  );
  X_BUF \_n0013<59>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<59>22_SW0/O ),
    .O(N5464)
  );
  defparam \_n0013<59>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<59>22_SW0  (
    .ADR0(data1[28]),
    .ADR1(_n0025),
    .ADR2(data1[60]),
    .ADR3(N01),
    .O(\_n0013<59>22_SW0/O )
  );
  X_BUF \_n0013<2>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<2>22_SW0/O ),
    .O(N5458)
  );
  defparam \_n0013<2>22_SW0 .INIT = 16'hEAC0;
  X_LUT4 \_n0013<2>22_SW0  (
    .ADR0(data1[3]),
    .ADR1(data1[17]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<2>22_SW0/O )
  );
  X_BUF \_n0013<62>14/LUT3_L_BUF  (
    .I(\_n0013<62>14/O ),
    .O(CHOICE32)
  );
  defparam \_n0013<62>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<62>14  (
    .ADR0(CHOICE30),
    .ADR1(data1[8]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<62>14/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<17>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<17>11_G/O ),
    .O(N5789)
  );
  defparam \c1/Mxor_OUTR_Result<17>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<17>11_G  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[50]),
    .ADR2(N5490),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_11 ),
    .O(\c1/Mxor_OUTR_Result<17>11_G/O )
  );
  X_BUF \_n0013<62>21/LUT3_L_BUF  (
    .I(\_n0013<62>21/O ),
    .O(_n0013[62])
  );
  defparam \_n0013<62>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<62>21  (
    .ADR0(CHOICE32),
    .ADR1(data1[63]),
    .ADR2(N01),
    .O(\_n0013<62>21/O )
  );
  X_BUF \_n0013<44>5/LUT4_L_BUF  (
    .I(\_n0013<44>5/O ),
    .O(CHOICE109)
  );
  defparam \_n0013<44>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<44>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[38]),
    .ADR2(state_FFd8),
    .ADR3(datain_45_IBUF),
    .O(\_n0013<44>5/O )
  );
  X_BUF \key2<2>961_G/LUT4_L_BUF  (
    .I(\key2<2>961_G/O ),
    .O(N5791)
  );
  defparam \key2<2>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<2>961_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out72 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out44 ),
    .O(\key2<2>961_G/O )
  );
  X_BUF \_n0013<60>5/LUT4_L_BUF  (
    .I(\_n0013<60>5/O ),
    .O(CHOICE37)
  );
  defparam \_n0013<60>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<60>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[34]),
    .ADR2(state_FFd8),
    .ADR3(datain_61_IBUF),
    .O(\_n0013<60>5/O )
  );
  X_BUF \key2<26>271_G/LUT4_L_BUF  (
    .I(\key2<26>271_G/O ),
    .O(N5793)
  );
  defparam \key2<26>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<26>271_G  (
    .ADR0(roundsel_3_8),
    .ADR1(\key1[16] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[15] ),
    .O(\key2<26>271_G/O )
  );
  X_BUF \_n0013<6>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<6>22_SW0/O ),
    .O(N5450)
  );
  defparam \_n0013<6>22_SW0 .INIT = 16'hEAC0;
  X_LUT4 \_n0013<6>22_SW0  (
    .ADR0(data1[7]),
    .ADR1(data1[1]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<6>22_SW0/O )
  );
  X_BUF \_n0013<44>14/LUT3_L_BUF  (
    .I(\_n0013<44>14/O ),
    .O(CHOICE113)
  );
  defparam \_n0013<44>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<44>14  (
    .ADR0(CHOICE111),
    .ADR1(data1[14]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<44>14/O )
  );
  X_BUF \key2<29>1181_G/LUT4_L_BUF  (
    .I(\key2<29>1181_G/O ),
    .O(N5795)
  );
  defparam \key2<29>1181_G .INIT = 16'h0E04;
  X_LUT4 \key2<29>1181_G  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out91 ),
    .ADR2(roundsel_3_14),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out23 ),
    .O(\key2<29>1181_G/O )
  );
  X_BUF \key2<15>12/LUT4_L_BUF  (
    .I(\key2<15>12/O ),
    .O(CHOICE585)
  );
  defparam \key2<15>12 .INIT = 16'hCA00;
  X_LUT4 \key2<15>12  (
    .ADR0(\key1[59] ),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_2_1),
    .O(\key2<15>12/O )
  );
  X_BUF \key2<15>1191_G/LUT4_L_BUF  (
    .I(\key2<15>1191_G/O ),
    .O(N5797)
  );
  defparam \key2<15>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<15>1191_G  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out26 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out65 ),
    .O(\key2<15>1191_G/O )
  );
  X_BUF \_n0013<60>14/LUT3_L_BUF  (
    .I(\_n0013<60>14/O ),
    .O(CHOICE41)
  );
  defparam \_n0013<60>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<60>14  (
    .ADR0(CHOICE39),
    .ADR1(data1[16]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<60>14/O )
  );
  X_BUF \_n0013<44>21/LUT3_L_BUF  (
    .I(\_n0013<44>21/O ),
    .O(_n0013[44])
  );
  defparam \_n0013<44>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<44>21  (
    .ADR0(CHOICE113),
    .ADR1(data1[45]),
    .ADR2(N01),
    .O(\_n0013<44>21/O )
  );
  X_BUF \key2<20>961_G/LUT4_L_BUF  (
    .I(\key2<20>961_G/O ),
    .O(N5799)
  );
  defparam \key2<20>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<20>961_G  (
    .ADR0(roundsel_3_13),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out47 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out49 ),
    .O(\key2<20>961_G/O )
  );
  X_BUF \_n0013<60>21/LUT3_L_BUF  (
    .I(\_n0013<60>21/O ),
    .O(_n0013[60])
  );
  defparam \_n0013<60>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<60>21  (
    .ADR0(CHOICE41),
    .ADR1(data1[61]),
    .ADR2(N01),
    .O(\_n0013<60>21/O )
  );
  X_BUF \key2<37>271_G/LUT4_L_BUF  (
    .I(\key2<37>271_G/O ),
    .O(N5801)
  );
  defparam \key2<37>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<37>271_G  (
    .ADR0(roundsel_33),
    .ADR1(\key1[21] ),
    .ADR2(roundsel_2_13),
    .ADR3(\key1[56] ),
    .O(\key2<37>271_G/O )
  );
  X_BUF \key2<11>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<11>110_SW01_G/O ),
    .O(N5803)
  );
  defparam \key2<11>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<11>110_SW01_G  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out46 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out66 ),
    .O(\key2<11>110_SW01_G/O )
  );
  X_BUF \key2<25>271_G/LUT4_L_BUF  (
    .I(\key2<25>271_G/O ),
    .O(N5805)
  );
  defparam \key2<25>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<25>271_G  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[22] ),
    .ADR2(roundsel_2_4),
    .ADR3(\key1[21] ),
    .O(\key2<25>271_G/O )
  );
  X_BUF \key2<11>961_G/LUT4_L_BUF  (
    .I(\key2<11>961_G/O ),
    .O(N5807)
  );
  defparam \key2<11>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<11>961_G  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out26 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out72 ),
    .O(\key2<11>961_G/O )
  );
  X_BUF \_n0013<58>5/LUT4_L_BUF  (
    .I(\_n0013<58>5/O ),
    .O(CHOICE46)
  );
  defparam \_n0013<58>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<58>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[18]),
    .ADR2(state_FFd8),
    .ADR3(datain_59_IBUF),
    .O(\_n0013<58>5/O )
  );
  X_BUF \_n0013<40>5/LUT4_L_BUF  (
    .I(\_n0013<40>5/O ),
    .O(CHOICE118)
  );
  defparam \_n0013<40>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<40>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[6]),
    .ADR2(state_FFd8),
    .ADR3(datain_41_IBUF),
    .O(\_n0013<40>5/O )
  );
  X_BUF \key2<39>90_SW01_G/LUT3_L_BUF  (
    .I(\key2<39>90_SW01_G/O ),
    .O(N5809)
  );
  defparam \key2<39>90_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<39>90_SW01_G  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out14 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out78 ),
    .O(\key2<39>90_SW01_G/O )
  );
  X_BUF \_n0013<61>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<61>22_SW0/O ),
    .O(N5462)
  );
  defparam \_n0013<61>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<61>22_SW0  (
    .ADR0(data1[30]),
    .ADR1(_n0025),
    .ADR2(data1[62]),
    .ADR3(N01),
    .O(\_n0013<61>22_SW0/O )
  );
  X_BUF \_n0013<51>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<51>22_SW0/O ),
    .O(N5468)
  );
  defparam \_n0013<51>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<51>22_SW0  (
    .ADR0(data1[20]),
    .ADR1(_n0025),
    .ADR2(data1[52]),
    .ADR3(N01),
    .O(\_n0013<51>22_SW0/O )
  );
  X_BUF \_n0013<58>14/LUT3_L_BUF  (
    .I(\_n0013<58>14/O ),
    .O(CHOICE50)
  );
  defparam \_n0013<58>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<58>14  (
    .ADR0(CHOICE48),
    .ADR1(data1[24]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<58>14/O )
  );
  X_BUF \_n0013<58>21/LUT3_L_BUF  (
    .I(\_n0013<58>21/O ),
    .O(_n0013[58])
  );
  defparam \_n0013<58>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<58>21  (
    .ADR0(CHOICE50),
    .ADR1(data1[59]),
    .ADR2(N01),
    .O(\_n0013<58>21/O )
  );
  X_BUF \_n0013<40>14/LUT3_L_BUF  (
    .I(\_n0013<40>14/O ),
    .O(CHOICE122)
  );
  defparam \_n0013<40>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<40>14  (
    .ADR0(CHOICE120),
    .ADR1(data1[30]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<40>14/O )
  );
  X_BUF \_n0013<0>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<0>22_SW0/O ),
    .O(N5456)
  );
  defparam \_n0013<0>22_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<0>22_SW0  (
    .ADR0(data1[25]),
    .ADR1(data1[1]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<0>22_SW0/O )
  );
  X_BUF \_n0013<40>21/LUT3_L_BUF  (
    .I(\_n0013<40>21/O ),
    .O(_n0013[40])
  );
  defparam \_n0013<40>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<40>21  (
    .ADR0(CHOICE122),
    .ADR1(data1[41]),
    .ADR2(N01),
    .O(\_n0013<40>21/O )
  );
  X_BUF \key2<23>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<23>133_SW01_G/O ),
    .O(N5811)
  );
  defparam \key2<23>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<23>133_SW01_G  (
    .ADR0(roundsel_2_8),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out35 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out34 ),
    .O(\key2<23>133_SW01_G/O )
  );
  X_BUF \key2<30>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<30>133_SW01_G/O ),
    .O(N5813)
  );
  defparam \key2<30>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<30>133_SW01_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out6 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out5 ),
    .O(\key2<30>133_SW01_G/O )
  );
  X_BUF \key2<46>1191_G/LUT4_L_BUF  (
    .I(\key2<46>1191_G/O ),
    .O(N5815)
  );
  defparam \key2<46>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<46>1191_G  (
    .ADR0(roundsel_3_14),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out84 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out86 ),
    .O(\key2<46>1191_G/O )
  );
  X_BUF \_n0013<54>5/LUT4_L_BUF  (
    .I(\_n0013<54>5/O ),
    .O(CHOICE55)
  );
  defparam \_n0013<54>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<54>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[52]),
    .ADR2(state_FFd8),
    .ADR3(datain_55_IBUF),
    .O(\_n0013<54>5/O )
  );
  X_BUF \_n0013<37>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<37>22_SW0/O ),
    .O(N5474)
  );
  defparam \_n0013<37>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<37>22_SW0  (
    .ADR0(data1[6]),
    .ADR1(_n0025),
    .ADR2(data1[38]),
    .ADR3(N01),
    .O(\_n0013<37>22_SW0/O )
  );
  X_BUF \key2<13>271_G/LUT4_L_BUF  (
    .I(\key2<13>271_G/O ),
    .O(N5817)
  );
  defparam \key2<13>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<13>271_G  (
    .ADR0(roundsel_3_6),
    .ADR1(\key1[3] ),
    .ADR2(roundsel_2_10),
    .ADR3(\key1[4] ),
    .O(\key2<13>271_G/O )
  );
  X_BUF \key2<42>961_G/LUT4_L_BUF  (
    .I(\key2<42>961_G/O ),
    .O(N5819)
  );
  defparam \key2<42>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<42>961_G  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out5 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out84 ),
    .O(\key2<42>961_G/O )
  );
  X_BUF \_n0013<38>5/LUT4_L_BUF  (
    .I(\_n0013<38>5/O ),
    .O(CHOICE127)
  );
  defparam \_n0013<38>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<38>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[56]),
    .ADR2(state_FFd8),
    .ADR3(datain_39_IBUF),
    .O(\_n0013<38>5/O )
  );
  X_BUF \_n0013<54>14/LUT3_L_BUF  (
    .I(\_n0013<54>14/O ),
    .O(CHOICE59)
  );
  defparam \_n0013<54>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<54>14  (
    .ADR0(CHOICE57),
    .ADR1(data1[7]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<54>14/O )
  );
  X_BUF \_n0013<9>20_SW0_SW0_SW0_SW0/LUT4_L_BUF  (
    .I(\_n0013<9>20_SW0_SW0_SW0_SW0/O ),
    .O(N5199)
  );
  defparam \_n0013<9>20_SW0_SW0_SW0_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<9>20_SW0_SW0_SW0_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1927),
    .ADR3(cipherout2[10]),
    .O(\_n0013<9>20_SW0_SW0_SW0_SW0/O )
  );
  X_BUF \key2<10>961_G/LUT4_L_BUF  (
    .I(\key2<10>961_G/O ),
    .O(N5821)
  );
  defparam \key2<10>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<10>961_G  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out33 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out47 ),
    .O(\key2<10>961_G/O )
  );
  X_BUF \_n0013<54>21/LUT3_L_BUF  (
    .I(\_n0013<54>21/O ),
    .O(_n0013[54])
  );
  defparam \_n0013<54>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<54>21  (
    .ADR0(CHOICE59),
    .ADR1(data1[55]),
    .ADR2(N01),
    .O(\_n0013<54>21/O )
  );
  X_BUF \key2<15>471_G/LUT4_L_BUF  (
    .I(\key2<15>471_G/O ),
    .O(N5823)
  );
  defparam \key2<15>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<15>471_G  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[42] ),
    .ADR2(roundsel_3_1),
    .ADR3(\key1[11] ),
    .O(\key2<15>471_G/O )
  );
  X_BUF \key2<9>1191_G/LUT4_L_BUF  (
    .I(\key2<9>1191_G/O ),
    .O(N5825)
  );
  defparam \key2<9>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<9>1191_G  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out28 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out66 ),
    .O(\key2<9>1191_G/O )
  );
  X_BUF \key2<27>471_G/LUT4_L_BUF  (
    .I(\key2<27>471_G/O ),
    .O(N5827)
  );
  defparam \key2<27>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<27>471_G  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[7] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[6] ),
    .O(\key2<27>471_G/O )
  );
  X_BUF \_n0013<38>14/LUT3_L_BUF  (
    .I(\_n0013<38>14/O ),
    .O(CHOICE131)
  );
  defparam \_n0013<38>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<38>14  (
    .ADR0(CHOICE129),
    .ADR1(data1[5]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<38>14/O )
  );
  X_BUF \_n0013<56>5/LUT4_L_BUF  (
    .I(\_n0013<56>5/O ),
    .O(CHOICE64)
  );
  defparam \_n0013<56>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<56>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[2]),
    .ADR2(state_FFd8),
    .ADR3(datain_57_IBUF),
    .O(\_n0013<56>5/O )
  );
  X_BUF \c1/Mxor_X_Result<31>11_G/LUT3_L_BUF  (
    .I(\c1/Mxor_X_Result<31>11_G/O ),
    .O(N5829)
  );
  defparam \c1/Mxor_X_Result<31>11_G .INIT = 8'h56;
  X_LUT3 \c1/Mxor_X_Result<31>11_G  (
    .ADR0(data1[12]),
    .ADR1(CHOICE1669),
    .ADR2(CHOICE1663),
    .O(\c1/Mxor_X_Result<31>11_G/O )
  );
  X_BUF \_n0013<39>12/LUT2_L_BUF  (
    .I(\_n0013<39>12/O ),
    .O(CHOICE788)
  );
  defparam \_n0013<39>12 .INIT = 4'h8;
  X_LUT2 \_n0013<39>12  (
    .ADR0(data1[40]),
    .ADR1(N01),
    .O(\_n0013<39>12/O )
  );
  X_BUF \_n0013<38>21/LUT3_L_BUF  (
    .I(\_n0013<38>21/O ),
    .O(_n0013[38])
  );
  defparam \_n0013<38>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<38>21  (
    .ADR0(CHOICE131),
    .ADR1(data1[39]),
    .ADR2(N01),
    .O(\_n0013<38>21/O )
  );
  X_BUF \key2<24>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<24>133_SW01_G/O ),
    .O(N5831)
  );
  defparam \key2<24>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<24>133_SW01_G  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out30 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out29 ),
    .O(\key2<24>133_SW01_G/O )
  );
  X_BUF \_n0013<56>14/LUT3_L_BUF  (
    .I(\_n0013<56>14/O ),
    .O(CHOICE68)
  );
  defparam \_n0013<56>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<56>14  (
    .ADR0(CHOICE66),
    .ADR1(data1[32]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<56>14/O )
  );
  X_BUF \key2<27>1411_G/LUT4_L_BUF  (
    .I(\key2<27>1411_G/O ),
    .O(N5833)
  );
  defparam \key2<27>1411_G .INIT = 16'h0E04;
  X_LUT4 \key2<27>1411_G  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out79 ),
    .O(\key2<27>1411_G/O )
  );
  X_BUF \key2<10>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<10>110_SW01_G/O ),
    .O(N5835)
  );
  defparam \key2<10>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<10>110_SW01_G  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out43 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out73 ),
    .O(\key2<10>110_SW01_G/O )
  );
  X_BUF \_n0013<56>21/LUT3_L_BUF  (
    .I(\_n0013<56>21/O ),
    .O(_n0013[56])
  );
  defparam \_n0013<56>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<56>21  (
    .ADR0(CHOICE68),
    .ADR1(data1[57]),
    .ADR2(N01),
    .O(\_n0013<56>21/O )
  );
  X_BUF \key2<2>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<2>110_SW01_G/O ),
    .O(N5837)
  );
  defparam \key2<2>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<2>110_SW01_G  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out54 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out61 ),
    .O(\key2<2>110_SW01_G/O )
  );
  X_BUF \key2<5>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<5>110_SW01_G/O ),
    .O(N5839)
  );
  defparam \key2<5>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<5>110_SW01_G  (
    .ADR0(roundsel_2_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out59 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .O(\key2<5>110_SW01_G/O )
  );
  X_BUF \_n0013<36>5/LUT4_L_BUF  (
    .I(\_n0013<36>5/O ),
    .O(CHOICE136)
  );
  defparam \_n0013<36>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<36>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[40]),
    .ADR2(state_FFd8),
    .ADR3(datain_37_IBUF),
    .O(\_n0013<36>5/O )
  );
  X_BUF \_n0013<10>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<10>22_SW0/O ),
    .O(N5454)
  );
  defparam \_n0013<10>22_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<10>22_SW0  (
    .ADR0(data1[18]),
    .ADR1(data1[11]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<10>22_SW0/O )
  );
  X_BUF \_n0013<18>17_SW0/LUT4_L_BUF  (
    .I(\_n0013<18>17_SW0/O ),
    .O(N5495)
  );
  defparam \_n0013<18>17_SW0 .INIT = 16'hFFA8;
  X_LUT4 \_n0013<18>17_SW0  (
    .ADR0(data1[19]),
    .ADR1(state_FFd7),
    .ADR2(N01),
    .ADR3(CHOICE616),
    .O(\_n0013<18>17_SW0/O )
  );
  X_BUF \_n0013<52>5/LUT4_L_BUF  (
    .I(\_n0013<52>5/O ),
    .O(CHOICE73)
  );
  defparam \_n0013<52>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<52>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[36]),
    .ADR2(state_FFd8),
    .ADR3(datain_53_IBUF),
    .O(\_n0013<52>5/O )
  );
  X_BUF \key2<7>761_G/LUT4_L_BUF  (
    .I(\key2<7>761_G/O ),
    .O(N5841)
  );
  defparam \key2<7>761_G .INIT = 16'h0E04;
  X_LUT4 \key2<7>761_G  (
    .ADR0(roundsel_33),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out65 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .O(\key2<7>761_G/O )
  );
  X_BUF \key2<33>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<33>110_SW01_G/O ),
    .O(N5843)
  );
  defparam \key2<33>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<33>110_SW01_G  (
    .ADR0(roundsel_3_2),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out22 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out86 ),
    .O(\key2<33>110_SW01_G/O )
  );
  X_BUF \key2<45>1191_G/LUT4_L_BUF  (
    .I(\key2<45>1191_G/O ),
    .O(N5845)
  );
  defparam \key2<45>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<45>1191_G  (
    .ADR0(roundsel_23),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out91 ),
    .ADR2(roundsel_3_14),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out84 ),
    .O(\key2<45>1191_G/O )
  );
  X_BUF \key2<5>961_G/LUT4_L_BUF  (
    .I(\key2<5>961_G/O ),
    .O(N5847)
  );
  defparam \key2<5>961_G .INIT = 16'h0E04;
  X_LUT4 \key2<5>961_G  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out39 ),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out41 ),
    .O(\key2<5>961_G/O )
  );
  X_BUF \key2<14>133_SW01_G/LUT3_L_BUF  (
    .I(\key2<14>133_SW01_G/O ),
    .O(N5849)
  );
  defparam \key2<14>133_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<14>133_SW01_G  (
    .ADR0(roundsel_3_13),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out36 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .O(\key2<14>133_SW01_G/O )
  );
  X_BUF \_n0013<36>14/LUT3_L_BUF  (
    .I(\_n0013<36>14/O ),
    .O(CHOICE140)
  );
  defparam \_n0013<36>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<36>14  (
    .ADR0(CHOICE138),
    .ADR1(data1[13]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<36>14/O )
  );
  X_BUF \_n0013<41>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<41>22_SW0/O ),
    .O(N5472)
  );
  defparam \_n0013<41>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<41>22_SW0  (
    .ADR0(data1[10]),
    .ADR1(_n0025),
    .ADR2(data1[42]),
    .ADR3(N01),
    .O(\_n0013<41>22_SW0/O )
  );
  X_BUF \_n0013<52>14/LUT3_L_BUF  (
    .I(\_n0013<52>14/O ),
    .O(CHOICE77)
  );
  defparam \_n0013<52>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<52>14  (
    .ADR0(CHOICE75),
    .ADR1(data1[15]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<52>14/O )
  );
  X_BUF \key2<43>271_G/LUT4_L_BUF  (
    .I(\key2<43>271_G/O ),
    .O(N5851)
  );
  defparam \key2<43>271_G .INIT = 16'h0E04;
  X_LUT4 \key2<43>271_G  (
    .ADR0(roundsel_3_6),
    .ADR1(\key1[46] ),
    .ADR2(roundsel_2_10),
    .ADR3(\key1[16] ),
    .O(\key2<43>271_G/O )
  );
  X_BUF \_n0013<55>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<55>22_SW0/O ),
    .O(N5466)
  );
  defparam \_n0013<55>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<55>22_SW0  (
    .ADR0(data1[24]),
    .ADR1(_n0025),
    .ADR2(data1[56]),
    .ADR3(N01),
    .O(\_n0013<55>22_SW0/O )
  );
  X_BUF \_n0013<36>21/LUT3_L_BUF  (
    .I(\_n0013<36>21/O ),
    .O(_n0013[36])
  );
  defparam \_n0013<36>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<36>21  (
    .ADR0(CHOICE140),
    .ADR1(data1[37]),
    .ADR2(N01),
    .O(\_n0013<36>21/O )
  );
  X_BUF \_n0013<52>21/LUT3_L_BUF  (
    .I(\_n0013<52>21/O ),
    .O(_n0013[52])
  );
  defparam \_n0013<52>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<52>21  (
    .ADR0(CHOICE77),
    .ADR1(data1[53]),
    .ADR2(N01),
    .O(\_n0013<52>21/O )
  );
  X_BUF \c1/Mxor_X_Result<15>11_G/LUT3_L_BUF  (
    .I(\c1/Mxor_X_Result<15>11_G/O ),
    .O(N5853)
  );
  defparam \c1/Mxor_X_Result<15>11_G .INIT = 8'h56;
  X_LUT3 \c1/Mxor_X_Result<15>11_G  (
    .ADR0(data1[22]),
    .ADR1(CHOICE503),
    .ADR2(CHOICE497),
    .O(\c1/Mxor_X_Result<15>11_G/O )
  );
  X_BUF \key2<28>471_G/LUT4_L_BUF  (
    .I(\key2<28>471_G/O ),
    .O(N5855)
  );
  defparam \key2<28>471_G .INIT = 16'h0E04;
  X_LUT4 \key2<28>471_G  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[7] ),
    .ADR2(roundsel_4_1),
    .ADR3(\key1[39] ),
    .O(\key2<28>471_G/O )
  );
  X_BUF \key2<17>1191_G/LUT4_L_BUF  (
    .I(\key2<17>1191_G/O ),
    .O(N5857)
  );
  defparam \key2<17>1191_G .INIT = 16'h0E04;
  X_LUT4 \key2<17>1191_G  (
    .ADR0(roundsel_2_8),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out61 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .O(\key2<17>1191_G/O )
  );
  X_BUF \key2<20>110_SW01_G/LUT3_L_BUF  (
    .I(\key2<20>110_SW01_G/O ),
    .O(N5859)
  );
  defparam \key2<20>110_SW01_G .INIT = 8'h27;
  X_LUT3 \key2<20>110_SW01_G  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out53 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out51 ),
    .O(\key2<20>110_SW01_G/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_291_G/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_291_G/O ),
    .O(N5861)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_291_G .INIT = 16'h3E94;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_291_G  (
    .ADR0(\c1/X[28] ),
    .ADR1(\c1/X[29] ),
    .ADR2(\c1/X[27] ),
    .ADR3(\c1/X[26] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_291_G/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_281_G/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_281_G/O ),
    .O(N5863)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_281_G .INIT = 16'h863D;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_281_G  (
    .ADR0(\c1/X[27] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[29] ),
    .ADR3(\c1/X[26] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_281_G/O )
  );
  X_BUF \_n0013<50>5/LUT4_L_BUF  (
    .I(\_n0013<50>5/O ),
    .O(CHOICE82)
  );
  defparam \_n0013<50>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<50>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[20]),
    .ADR2(state_FFd8),
    .ADR3(datain_51_IBUF),
    .O(\_n0013<50>5/O )
  );
  X_BUF \_n0013<32>5/LUT4_L_BUF  (
    .I(\_n0013<32>5/O ),
    .O(CHOICE145)
  );
  defparam \_n0013<32>5 .INIT = 16'hF888;
  X_LUT4 \_n0013<32>5  (
    .ADR0(state_FFd7),
    .ADR1(data1[8]),
    .ADR2(state_FFd8),
    .ADR3(datain_33_IBUF),
    .O(\_n0013<32>5/O )
  );
  X_BUF \roundsel<2>_mmx_out331_G/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out331_G/O ),
    .O(N5865)
  );
  defparam \roundsel<2>_mmx_out331_G .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out331_G  (
    .ADR0(roundsel_1_11),
    .ADR1(\key1[59] ),
    .ADR2(\key1[12] ),
    .O(\roundsel<2>_mmx_out331_G/O )
  );
  X_BUF \_n0013<50>14/LUT3_L_BUF  (
    .I(\_n0013<50>14/O ),
    .O(CHOICE86)
  );
  defparam \_n0013<50>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<50>14  (
    .ADR0(CHOICE84),
    .ADR1(data1[23]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<50>14/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_251_G/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_251_G/O ),
    .O(N5867)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_251_G .INIT = 16'hEA25;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_251_G  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[29] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_251_G/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_241_G/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_241_G/O ),
    .O(N5869)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_241_G .INIT = 16'h26BC;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_241_G  (
    .ADR0(\c1/X[28] ),
    .ADR1(\c1/X[29] ),
    .ADR2(\c1/X[26] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_241_G/O )
  );
  X_BUF \_n0013<50>21/LUT3_L_BUF  (
    .I(\_n0013<50>21/O ),
    .O(_n0013[50])
  );
  defparam \_n0013<50>21 .INIT = 8'hEA;
  X_LUT3 \_n0013<50>21  (
    .ADR0(CHOICE86),
    .ADR1(data1[51]),
    .ADR2(N01),
    .O(\_n0013<50>21/O )
  );
  X_BUF \c1/u6/Mrom_dout_inst_mux_f5_111_G/LUT4_L_BUF  (
    .I(\c1/u6/Mrom_dout_inst_mux_f5_111_G/O ),
    .O(N5871)
  );
  defparam \c1/u6/Mrom_dout_inst_mux_f5_111_G .INIT = 16'h69C9;
  X_LUT4 \c1/u6/Mrom_dout_inst_mux_f5_111_G  (
    .ADR0(\c1/X[39] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[38] ),
    .O(\c1/u6/Mrom_dout_inst_mux_f5_111_G/O )
  );
  X_BUF \_n0013<32>14/LUT3_L_BUF  (
    .I(\_n0013<32>14/O ),
    .O(CHOICE149)
  );
  defparam \_n0013<32>14 .INIT = 8'hEA;
  X_LUT3 \_n0013<32>14  (
    .ADR0(CHOICE147),
    .ADR1(data1[29]),
    .ADR2(\state_FFd3-In ),
    .O(\_n0013<32>14/O )
  );
  X_BUF \Ker020_SW0/LUT3_L_BUF  (
    .I(\Ker020_SW0/O ),
    .O(N5428)
  );
  defparam Ker020_SW0.INIT = 8'hFE;
  X_LUT3 Ker020_SW0 (
    .ADR0(state_FFd2),
    .ADR1(state_FFd6),
    .ADR2(state_FFd4),
    .O(\Ker020_SW0/O )
  );
  X_BUF \_n0013<26>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<26>22_SW0/O ),
    .O(N5478)
  );
  defparam \_n0013<26>22_SW0 .INIT = 16'hEAC0;
  X_LUT4 \_n0013<26>22_SW0  (
    .ADR0(data1[27]),
    .ADR1(data1[20]),
    .ADR2(\state_FFd3-In ),
    .ADR3(N01),
    .O(\_n0013<26>22_SW0/O )
  );
  X_BUF \_n0013<7>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<7>20_SW0/O ),
    .O(N5430)
  );
  defparam \_n0013<7>20_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<7>20_SW0  (
    .ADR0(data1[8]),
    .ADR1(_n0025),
    .ADR2(N01),
    .ADR3(cipherout2[8]),
    .O(\_n0013<7>20_SW0/O )
  );
  X_BUF \c1/u6/Mrom_dout_inst_mux_f5_101_G/LUT4_L_BUF  (
    .I(\c1/u6/Mrom_dout_inst_mux_f5_101_G/O ),
    .O(N5873)
  );
  defparam \c1/u6/Mrom_dout_inst_mux_f5_101_G .INIT = 16'hE466;
  X_LUT4 \c1/u6/Mrom_dout_inst_mux_f5_101_G  (
    .ADR0(\c1/X[39] ),
    .ADR1(\c1/X[41] ),
    .ADR2(\c1/X[38] ),
    .ADR3(\c1/X[40] ),
    .O(\c1/u6/Mrom_dout_inst_mux_f5_101_G/O )
  );
  X_BUF \_n0013<15>20/LUT4_L_BUF  (
    .I(\_n0013<15>20/O ),
    .O(_n0013[15])
  );
  defparam \_n0013<15>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<15>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE2009),
    .ADR2(cipherout2[2]),
    .ADR3(N5039),
    .O(\_n0013<15>20/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<25>11_G/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<25>11_G/O ),
    .O(N5875)
  );
  defparam \c1/Mxor_OUTR_Result<25>11_G .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<25>11_G  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[58]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_29 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_31 ),
    .O(\c1/Mxor_OUTR_Result<25>11_G/O )
  );
  X_BUF \_n0013<27>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<27>20_SW0/O ),
    .O(N5019)
  );
  defparam \_n0013<27>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<27>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1972),
    .ADR3(cipherout2[28]),
    .O(\_n0013<27>20_SW0/O )
  );
  X_BUF \roundsel<2>_mmx_out241_G/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out241_G/O ),
    .O(N5877)
  );
  defparam \roundsel<2>_mmx_out241_G .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out241_G  (
    .ADR0(roundsel_11),
    .ADR1(\key1[12] ),
    .ADR2(\key1[28] ),
    .O(\roundsel<2>_mmx_out241_G/O )
  );
  X_BUF \key2<31>15_G/LUT4_L_BUF  (
    .I(\key2<31>15_G/O ),
    .O(N5879)
  );
  defparam \key2<31>15_G .INIT = 16'h0E04;
  X_LUT4 \key2<31>15_G  (
    .ADR0(roundsel_1_7),
    .ADR1(\key1[21] ),
    .ADR2(roundsel_3_16),
    .ADR3(\key1[8] ),
    .O(\key2<31>15_G/O )
  );
  X_BUF \key2<9>12/LUT4_L_BUF  (
    .I(\key2<9>12/O ),
    .O(CHOICE1411)
  );
  defparam \key2<9>12 .INIT = 16'hAC00;
  X_LUT4 \key2<9>12  (
    .ADR0(\key1[61] ),
    .ADR1(\key1[53] ),
    .ADR2(roundsel_1_10),
    .ADR3(roundsel_3_5),
    .O(\key2<9>12/O )
  );
  X_BUF \_n0013<3>20/LUT4_L_BUF  (
    .I(\_n0013<3>20/O ),
    .O(_n0013[3])
  );
  defparam \_n0013<3>20 .INIT = 16'hFFEA;
  X_LUT4 \_n0013<3>20  (
    .ADR0(CHOICE1345),
    .ADR1(_n0025),
    .ADR2(cipherout2[4]),
    .ADR3(N5434),
    .O(\_n0013<3>20/O )
  );
  X_BUF \key2<46>12/LUT4_L_BUF  (
    .I(\key2<46>12/O ),
    .O(CHOICE1887)
  );
  defparam \key2<46>12 .INIT = 16'hCA00;
  X_LUT4 \key2<46>12  (
    .ADR0(\key1[15] ),
    .ADR1(\key1[23] ),
    .ADR2(roundsel_1_6),
    .ADR3(roundsel_3_1),
    .O(\key2<46>12/O )
  );
  X_BUF \key2<26>12_G/LUT4_L_BUF  (
    .I(\key2<26>12_G/O ),
    .O(N5881)
  );
  defparam \key2<26>12_G .INIT = 16'hA280;
  X_LUT4 \key2<26>12_G  (
    .ADR0(roundsel_2_6),
    .ADR1(roundsel_1_18),
    .ADR2(\key1[39] ),
    .ADR3(\key1[31] ),
    .O(\key2<26>12_G/O )
  );
  X_BUF \_n0013<11>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<11>20_SW0/O ),
    .O(N5047)
  );
  defparam \_n0013<11>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<11>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1936),
    .ADR3(cipherout2[12]),
    .O(\_n0013<11>20_SW0/O )
  );
  X_BUF \_n0013<1>20/LUT4_L_BUF  (
    .I(\_n0013<1>20/O ),
    .O(_n0013[1])
  );
  defparam \_n0013<1>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<1>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1946),
    .ADR2(cipherout2[25]),
    .ADR3(N5033),
    .O(\_n0013<1>20/O )
  );
  X_BUF \_n0013<19>20/LUT4_L_BUF  (
    .I(\_n0013<19>20/O ),
    .O(_n0013[19])
  );
  defparam \_n0013<19>20 .INIT = 16'hFFEA;
  X_LUT4 \_n0013<19>20  (
    .ADR0(CHOICE1999),
    .ADR1(_n0025),
    .ADR2(cipherout2[20]),
    .ADR3(N5436),
    .O(\_n0013<19>20/O )
  );
  X_BUF \key2<19>12/LUT4_D_BUF  (
    .I(CHOICE849),
    .O(N5940)
  );
  defparam \key2<19>12 .INIT = 16'hA280;
  X_LUT4 \key2<19>12  (
    .ADR0(roundsel[3]),
    .ADR1(roundsel[2]),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out56 ),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out39 ),
    .O(CHOICE849)
  );
  X_BUF \_n0013<9>20/LUT4_L_BUF  (
    .I(\_n0013<9>20/O ),
    .O(_n0013[9])
  );
  defparam \_n0013<9>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<9>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1928),
    .ADR2(cipherout2[26]),
    .ADR3(N5199),
    .O(\_n0013<9>20/O )
  );
  X_BUF \_n0013<19>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<19>20_SW0/O ),
    .O(N5436)
  );
  defparam \_n0013<19>20_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<19>20_SW0  (
    .ADR0(data1[20]),
    .ADR1(\state_FFd3-In ),
    .ADR2(N01),
    .ADR3(cipherout2[19]),
    .O(\_n0013<19>20_SW0/O )
  );
  X_BUF \key2<8>12_G/LUT4_L_BUF  (
    .I(\key2<8>12_G/O ),
    .O(N5883)
  );
  defparam \key2<8>12_G .INIT = 16'hA280;
  X_LUT4 \key2<8>12_G  (
    .ADR0(roundsel_2_8),
    .ADR1(roundsel_1_5),
    .ADR2(\key1[42] ),
    .ADR3(\key1[34] ),
    .O(\key2<8>12_G/O )
  );
  X_BUF \_n0013<21>20/LUT4_L_BUF  (
    .I(\_n0013<21>20/O ),
    .O(_n0013[21])
  );
  defparam \_n0013<21>20 .INIT = 16'hFFEA;
  X_LUT4 \_n0013<21>20  (
    .ADR0(CHOICE1990),
    .ADR1(_n0025),
    .ADR2(cipherout2[22]),
    .ADR3(N5438),
    .O(\_n0013<21>20/O )
  );
  X_BUF \_n0013<21>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<21>20_SW0/O ),
    .O(N5438)
  );
  defparam \_n0013<21>20_SW0 .INIT = 16'hECA0;
  X_LUT4 \_n0013<21>20_SW0  (
    .ADR0(data1[22]),
    .ADR1(\state_FFd3-In ),
    .ADR2(N01),
    .ADR3(cipherout2[11]),
    .O(\_n0013<21>20_SW0/O )
  );
  X_BUF \_n0013<23>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<23>20_SW0/O ),
    .O(N5035)
  );
  defparam \_n0013<23>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<23>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1276),
    .ADR3(cipherout2[24]),
    .O(\_n0013<23>20_SW0/O )
  );
  X_BUF \_n0013<25>20/LUT4_L_BUF  (
    .I(\_n0013<25>20/O ),
    .O(_n0013[25])
  );
  defparam \_n0013<25>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<25>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1982),
    .ADR2(cipherout2[28]),
    .ADR3(N5045),
    .O(\_n0013<25>20/O )
  );
  X_BUF \key2<37>12_SW0_G/LUT3_L_BUF  (
    .I(\key2<37>12_SW0_G/O ),
    .O(N5885)
  );
  defparam \key2<37>12_SW0_G .INIT = 8'hE4;
  X_LUT3 \key2<37>12_SW0_G  (
    .ADR0(roundsel_1_14),
    .ADR1(\key1[7] ),
    .ADR2(\key1[15] ),
    .O(\key2<37>12_SW0_G/O )
  );
  X_BUF \_n0013<15>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<15>20_SW0/O ),
    .O(N5039)
  );
  defparam \_n0013<15>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<15>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE2008),
    .ADR3(cipherout2[16]),
    .O(\_n0013<15>20_SW0/O )
  );
  X_BUF \_n0013<29>20/LUT4_L_BUF  (
    .I(\_n0013<29>20/O ),
    .O(_n0013[29])
  );
  defparam \_n0013<29>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<29>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1955),
    .ADR2(cipherout2[12]),
    .ADR3(N5151),
    .O(\_n0013<29>20/O )
  );
  X_BUF \_n0013<20>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<20>22_SW0/O ),
    .O(N5484)
  );
  defparam \_n0013<20>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<20>22_SW0  (
    .ADR0(data1[11]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[21]),
    .ADR3(N01),
    .O(\_n0013<20>22_SW0/O )
  );
  X_BUF \_n0013<16>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<16>22_SW0/O ),
    .O(N5486)
  );
  defparam \_n0013<16>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<16>22_SW0  (
    .ADR0(data1[27]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[17]),
    .ADR3(N01),
    .O(\_n0013<16>22_SW0/O )
  );
  X_BUF \_n0013<17>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<17>20_SW0/O ),
    .O(N5017)
  );
  defparam \_n0013<17>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<17>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1046),
    .ADR3(cipherout2[18]),
    .O(\_n0013<17>20_SW0/O )
  );
  X_BUF \_n0013<5>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<5>20_SW0/O ),
    .O(N5021)
  );
  defparam \_n0013<5>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<5>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1267),
    .ADR3(cipherout2[6]),
    .O(\_n0013<5>20_SW0/O )
  );
  X_BUF \_n0013<27>20/LUT4_L_BUF  (
    .I(\_n0013<27>20/O ),
    .O(_n0013[27])
  );
  defparam \_n0013<27>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<27>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1973),
    .ADR2(cipherout2[20]),
    .ADR3(N5019),
    .O(\_n0013<27>20/O )
  );
  X_BUF \key2<43>12_SW0_G/LUT3_L_BUF  (
    .I(\key2<43>12_SW0_G/O ),
    .O(N5887)
  );
  defparam \key2<43>12_SW0_G .INIT = 8'hE4;
  X_LUT3 \key2<43>12_SW0_G  (
    .ADR0(roundsel_1_14),
    .ADR1(\key1[32] ),
    .ADR2(\key1[40] ),
    .O(\key2<43>12_SW0_G/O )
  );
  X_BUF \_n0013<25>20_SW0/LUT4_L_BUF  (
    .I(\_n0013<25>20_SW0/O ),
    .O(N5045)
  );
  defparam \_n0013<25>20_SW0 .INIT = 16'hFEF0;
  X_LUT4 \_n0013<25>20_SW0  (
    .ADR0(state_FFd5),
    .ADR1(state_FFd6),
    .ADR2(CHOICE1981),
    .ADR3(cipherout2[26]),
    .O(\_n0013<25>20_SW0/O )
  );
  X_BUF \_n0013<5>20/LUT4_L_BUF  (
    .I(\_n0013<5>20/O ),
    .O(_n0013[5])
  );
  defparam \_n0013<5>20 .INIT = 16'hFFEC;
  X_LUT4 \_n0013<5>20  (
    .ADR0(\state_FFd3-In ),
    .ADR1(CHOICE1268),
    .ADR2(cipherout2[9]),
    .ADR3(N5021),
    .O(\_n0013<5>20/O )
  );
  X_BUF \_n0013<12>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<12>22_SW0/O ),
    .O(N5488)
  );
  defparam \_n0013<12>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<12>22_SW0  (
    .ADR0(data1[10]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[13]),
    .ADR3(N01),
    .O(\_n0013<12>22_SW0/O )
  );
  X_BUF \key2<13>12_SW0_G/LUT3_L_BUF  (
    .I(\key2<13>12_SW0_G/O ),
    .O(N5889)
  );
  defparam \key2<13>12_SW0_G .INIT = 8'hE4;
  X_LUT3 \key2<13>12_SW0_G  (
    .ADR0(roundsel_1_14),
    .ADR1(\key1[20] ),
    .ADR2(\key1[28] ),
    .O(\key2<13>12_SW0_G/O )
  );
  X_BUF \_n0013<22>22_SW0/LUT4_L_BUF  (
    .I(\_n0013<22>22_SW0/O ),
    .O(N5482)
  );
  defparam \_n0013<22>22_SW0 .INIT = 16'hF888;
  X_LUT4 \_n0013<22>22_SW0  (
    .ADR0(data1[3]),
    .ADR1(\state_FFd3-In ),
    .ADR2(data1[23]),
    .ADR3(N01),
    .O(\_n0013<22>22_SW0/O )
  );
  X_BUF \_n0013<31>20/LUT4_L_BUF  (
    .I(\_n0013<31>20/O ),
    .O(_n0013[31])
  );
  defparam \_n0013<31>20 .INIT = 16'hFAF8;
  X_LUT4 \_n0013<31>20  (
    .ADR0(cipherout2[32]),
    .ADR1(state_FFd5),
    .ADR2(N5193),
    .ADR3(state_FFd6),
    .O(\_n0013<31>20/O )
  );
  X_BUF \Ker039_1/LUT4_L_BUF  (
    .I(\Ker039_1/O ),
    .O(Ker039)
  );
  defparam Ker039_1.INIT = 16'hFFF2;
  X_LUT4 Ker039_1 (
    .ADR0(state_FFd2),
    .ADR1(_n0001),
    .ADR2(CHOICE195),
    .ADR3(CHOICE199),
    .O(\Ker039_1/O )
  );
  X_BUF \key2<7>15_G/LUT4_L_BUF  (
    .I(\key2<7>15_G/O ),
    .O(N5891)
  );
  defparam \key2<7>15_G .INIT = 16'h0E04;
  X_LUT4 \key2<7>15_G  (
    .ADR0(roundsel_11),
    .ADR1(\key1[59] ),
    .ADR2(roundsel_3_6),
    .ADR3(\key1[12] ),
    .O(\key2<7>15_G/O )
  );
  X_BUF \key2<26>61_G/LUT3_L_BUF  (
    .I(\key2<26>61_G/O ),
    .O(N5893)
  );
  defparam \key2<26>61_G .INIT = 8'hE4;
  X_LUT3 \key2<26>61_G  (
    .ADR0(roundsel_1_1),
    .ADR1(\key1[6] ),
    .ADR2(\key1[22] ),
    .O(\key2<26>61_G/O )
  );
  X_BUF \key2<31>12_G/LUT4_L_BUF  (
    .I(\key2<31>12_G/O ),
    .O(N5895)
  );
  defparam \key2<31>12_G .INIT = 16'hA280;
  X_LUT4 \key2<31>12_G  (
    .ADR0(roundsel_3_6),
    .ADR1(roundsel_1_4),
    .ADR2(\key1[64] ),
    .ADR3(\key1[56] ),
    .O(\key2<31>12_G/O )
  );
  X_BUF \key2<7>12_G/LUT4_L_BUF  (
    .I(\key2<7>12_G/O ),
    .O(N5897)
  );
  defparam \key2<7>12_G .INIT = 16'hA280;
  X_LUT4 \key2<7>12_G  (
    .ADR0(roundsel_3_6),
    .ADR1(roundsel_1_15),
    .ADR2(\key1[37] ),
    .ADR3(\key1[60] ),
    .O(\key2<7>12_G/O )
  );
  X_BUF \key2<22>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<22>110_SW01_F/O ),
    .O(N5620)
  );
  defparam \key2<22>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<22>110_SW01_F  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out41 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out38 ),
    .O(\key2<22>110_SW01_F/O )
  );
  X_BUF \key2<4>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<4>110_SW01_F/O ),
    .O(N5622)
  );
  defparam \key2<4>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<4>110_SW01_F  (
    .ADR0(roundsel_3_5),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out24 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .O(\key2<4>110_SW01_F/O )
  );
  X_BUF \key2<3>1181_F/LUT4_L_BUF  (
    .I(\key2<3>1181_F/O ),
    .O(N5624)
  );
  defparam \key2<3>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<3>1181_F  (
    .ADR0(roundsel_4_6),
    .ADR1(CHOICE1577),
    .ADR2(roundsel_2_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out47 ),
    .O(\key2<3>1181_F/O )
  );
  X_BUF \key2<32>271_F/LUT4_L_BUF  (
    .I(\key2<32>271_F/O ),
    .O(N5626)
  );
  defparam \key2<32>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<32>271_F  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[39] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[38] ),
    .O(\key2<32>271_F/O )
  );
  X_BUF \key2<47>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<47>110_SW01_F/O ),
    .O(N5628)
  );
  defparam \key2<47>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<47>110_SW01_F  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out81 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out79 ),
    .O(\key2<47>110_SW01_F/O )
  );
  X_BUF \key2<28>1191_F/LUT4_L_BUF  (
    .I(\key2<28>1191_F/O ),
    .O(N5630)
  );
  defparam \key2<28>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<28>1191_F  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out1 ),
    .ADR2(roundsel_3_15),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out20 ),
    .O(\key2<28>1191_F/O )
  );
  X_BUF \key2<25>961_F/LUT4_L_BUF  (
    .I(\key2<25>961_F/O ),
    .O(N5634)
  );
  defparam \key2<25>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<25>961_F  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out22 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out10 ),
    .O(\key2<25>961_F/O )
  );
  X_BUF \key2<37>961_F/LUT4_L_BUF  (
    .I(\key2<37>961_F/O ),
    .O(N5636)
  );
  defparam \key2<37>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<37>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out18 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .O(\key2<37>961_F/O )
  );
  X_BUF \key2<38>961_F/LUT4_L_BUF  (
    .I(\key2<38>961_F/O ),
    .O(N5638)
  );
  defparam \key2<38>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<38>961_F  (
    .ADR0(roundsel_3_5),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out16 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out31 ),
    .O(\key2<38>961_F/O )
  );
  X_BUF \key2<3>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<3>133_SW01_F/O ),
    .O(N5640)
  );
  defparam \key2<3>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<3>133_SW01_F  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out48 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out66 ),
    .O(\key2<3>133_SW01_F/O )
  );
  X_BUF \key2<25>12_SW0_F/LUT3_L_BUF  (
    .I(\key2<25>12_SW0_F/O ),
    .O(N5642)
  );
  defparam \key2<25>12_SW0_F .INIT = 8'hE4;
  X_LUT3 \key2<25>12_SW0_F  (
    .ADR0(roundsel_1_8),
    .ADR1(\key1[38] ),
    .ADR2(\key1[54] ),
    .O(\key2<25>12_SW0_F/O )
  );
  X_BUF \key2<21>1191_F/LUT4_L_BUF  (
    .I(\key2<21>1191_F/O ),
    .O(N5644)
  );
  defparam \key2<21>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<21>1191_F  (
    .ADR0(roundsel_2_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out43 ),
    .ADR2(roundsel_3_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out44 ),
    .O(\key2<21>1191_F/O )
  );
  X_BUF \key2<33>961_F/LUT4_L_BUF  (
    .I(\key2<33>961_F/O ),
    .O(N5646)
  );
  defparam \key2<33>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<33>961_F  (
    .ADR0(roundsel_3_2),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out14 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out81 ),
    .O(\key2<33>961_F/O )
  );
  X_BUF \roundsel<2>_mmx_out271_F/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out271_F/O ),
    .O(N5648)
  );
  defparam \roundsel<2>_mmx_out271_F .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out271_F  (
    .ADR0(roundsel_11),
    .ADR1(\key1[18] ),
    .ADR2(\key1[34] ),
    .O(\roundsel<2>_mmx_out271_F/O )
  );
  X_BUF \key2<22>961_F/LUT4_L_BUF  (
    .I(\key2<22>961_F/O ),
    .O(N5650)
  );
  defparam \key2<22>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<22>961_F  (
    .ADR0(roundsel_3_13),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out36 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out32 ),
    .O(\key2<22>961_F/O )
  );
  X_BUF \key2<32>12_F/LUT4_L_BUF  (
    .I(\key2<32>12_F/O ),
    .O(N5652)
  );
  defparam \key2<32>12_F .INIT = 16'hA280;
  X_LUT4 \key2<32>12_F  (
    .ADR0(roundsel_2_4),
    .ADR1(roundsel_1_20),
    .ADR2(\key1[22] ),
    .ADR3(\key1[6] ),
    .O(\key2<32>12_F/O )
  );
  X_BUF \roundsel<2>_mmx_out71_F/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out71_F/O ),
    .O(N5654)
  );
  defparam \roundsel<2>_mmx_out71_F .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out71_F  (
    .ADR0(roundsel_1_8),
    .ADR1(\key1[38] ),
    .ADR2(\key1[54] ),
    .O(\roundsel<2>_mmx_out71_F/O )
  );
  X_BUF \key2<29>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<29>133_SW01_F/O ),
    .O(N5656)
  );
  defparam \key2<29>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<29>133_SW01_F  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out87 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out84 ),
    .O(\key2<29>133_SW01_F/O )
  );
  X_BUF \key2<41>961_F/LUT4_L_BUF  (
    .I(\key2<41>961_F/O ),
    .O(N5658)
  );
  defparam \key2<41>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<41>961_F  (
    .ADR0(roundsel_3_10),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out7 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out80 ),
    .O(\key2<41>961_F/O )
  );
  X_BUF \key2<19>761_F/LUT4_L_BUF  (
    .I(\key2<19>761_F/O ),
    .O(N5660)
  );
  defparam \key2<19>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<19>761_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out54 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out37 ),
    .O(\key2<19>761_F/O )
  );
  X_BUF \roundsel<2>_mmx_out111_F/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out111_F/O ),
    .O(N5662)
  );
  defparam \roundsel<2>_mmx_out111_F .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out111_F  (
    .ADR0(roundsel_1_7),
    .ADR1(\key1[48] ),
    .ADR2(\key1[64] ),
    .O(\roundsel<2>_mmx_out111_F/O )
  );
  X_BUF \key2<39>761_F/LUT4_L_BUF  (
    .I(\key2<39>761_F/O ),
    .O(N5664)
  );
  defparam \key2<39>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<39>761_F  (
    .ADR0(roundsel_3_14),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out12 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .O(\key2<39>761_F/O )
  );
  X_BUF \key2<31>761_F/LUT4_L_BUF  (
    .I(\key2<31>761_F/O ),
    .O(N5666)
  );
  defparam \key2<31>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<31>761_F  (
    .ADR0(roundsel_3_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out19 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out94 ),
    .O(\key2<31>761_F/O )
  );
  X_BUF \key2<4>961_F/LUT4_L_BUF  (
    .I(\key2<4>961_F/O ),
    .O(N5668)
  );
  defparam \key2<4>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<4>961_F  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out35 ),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out73 ),
    .O(\key2<4>961_F/O )
  );
  X_BUF \key2<47>961_F/LUT4_L_BUF  (
    .I(\key2<47>961_F/O ),
    .O(N5670)
  );
  defparam \key2<47>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<47>961_F  (
    .ADR0(roundsel_3_5),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out76 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out78 ),
    .O(\key2<47>961_F/O )
  );
  X_BUF \key2<44>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<44>110_SW01_F/O ),
    .O(N5672)
  );
  defparam \key2<44>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<44>110_SW01_F  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out94 ),
    .O(\key2<44>110_SW01_F/O )
  );
  X_BUF \key2<34>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<34>110_SW01_F/O ),
    .O(N5674)
  );
  defparam \key2<34>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<34>110_SW01_F  (
    .ADR0(roundsel_3_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out5 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out9 ),
    .O(\key2<34>110_SW01_F/O )
  );
  X_BUF \key2<43>961_F/LUT4_L_BUF  (
    .I(\key2<43>961_F/O ),
    .O(N5676)
  );
  defparam \key2<43>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<43>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out2 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out93 ),
    .O(\key2<43>961_F/O )
  );
  X_BUF \c1/Mxor_X_Result<7>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_X_Result<7>11_F/O ),
    .O(N5678)
  );
  defparam \c1/Mxor_X_Result<7>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_X_Result<7>11_F  (
    .ADR0(roundsel[3]),
    .ADR1(data1[28]),
    .ADR2(CHOICE1628),
    .ADR3(\MUX_BLOCK_roundsel<2>_mmx_out24 ),
    .O(\c1/Mxor_X_Result<7>11_F/O )
  );
  X_BUF \key2<35>761_F/LUT4_L_BUF  (
    .I(\key2<35>761_F/O ),
    .O(N5680)
  );
  defparam \key2<35>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<35>761_F  (
    .ADR0(roundsel_3_2),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out17 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out9 ),
    .O(\key2<35>761_F/O )
  );
  X_BUF \key2<45>471_F/LUT4_L_BUF  (
    .I(\key2<45>471_F/O ),
    .O(N5682)
  );
  defparam \key2<45>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<45>471_F  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[32] ),
    .ADR2(roundsel_4_1),
    .ADR3(\key1[64] ),
    .O(\key2<45>471_F/O )
  );
  X_BUF \key2<6>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<6>110_SW01_F/O ),
    .O(N5684)
  );
  defparam \key2<6>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<6>110_SW01_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out44 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out72 ),
    .O(\key2<6>110_SW01_F/O )
  );
  X_BUF \key2<34>961_F/LUT4_L_BUF  (
    .I(\key2<34>961_F/O ),
    .O(N5686)
  );
  defparam \key2<34>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<34>961_F  (
    .ADR0(roundsel_3_8),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out64 ),
    .ADR2(roundsel_4_2),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out95 ),
    .O(\key2<34>961_F/O )
  );
  X_BUF \key2<6>961_F/LUT4_L_BUF  (
    .I(\key2<6>961_F/O ),
    .O(N5688)
  );
  defparam \key2<6>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<6>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out69 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out41 ),
    .O(\key2<6>961_F/O )
  );
  X_BUF \key2<35>90_SW01_F/LUT3_L_BUF  (
    .I(\key2<35>90_SW01_F/O ),
    .O(N5690)
  );
  defparam \key2<35>90_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<35>90_SW01_F  (
    .ADR0(roundsel_3_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out88 ),
    .O(\key2<35>90_SW01_F/O )
  );
  X_BUF \key2<30>1181_F/LUT4_L_BUF  (
    .I(\key2<30>1181_F/O ),
    .O(N5692)
  );
  defparam \key2<30>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<30>1181_F  (
    .ADR0(roundsel[3]),
    .ADR1(CHOICE455),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out ),
    .O(\key2<30>1181_F/O )
  );
  X_BUF \key2<17>471_F/LUT4_L_BUF  (
    .I(\key2<17>471_F/O ),
    .O(N5694)
  );
  defparam \key2<17>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<17>471_F  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[53] ),
    .ADR2(roundsel_3_1),
    .ADR3(\key1[18] ),
    .O(\key2<17>471_F/O )
  );
  X_BUF \key2<18>961_F/LUT4_L_BUF  (
    .I(\key2<18>961_F/O ),
    .O(N5696)
  );
  defparam \key2<18>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<18>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out57 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out51 ),
    .O(\key2<18>961_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<16>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<16>11_F/O ),
    .O(N5698)
  );
  defparam \c1/Mxor_OUTR_Result<16>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<16>11_F  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[49]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_84 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_86 ),
    .O(\c1/Mxor_OUTR_Result<16>11_F/O )
  );
  X_BUF \key2<42>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<42>110_SW01_F/O ),
    .O(N5700)
  );
  defparam \key2<42>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<42>110_SW01_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out23 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out15 ),
    .O(\key2<42>110_SW01_F/O )
  );
  X_BUF \key2<40>90_SW01_F/LUT3_L_BUF  (
    .I(\key2<40>90_SW01_F/O ),
    .O(N5702)
  );
  defparam \key2<40>90_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<40>90_SW01_F  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out10 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out86 ),
    .O(\key2<40>90_SW01_F/O )
  );
  X_BUF \key2<21>471_F/LUT4_L_BUF  (
    .I(\key2<21>471_F/O ),
    .O(N5704)
  );
  defparam \key2<21>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<21>471_F  (
    .ADR0(roundsel_2_4),
    .ADR1(\key1[4] ),
    .ADR2(roundsel_4_2),
    .ADR3(\key1[36] ),
    .O(\key2<21>471_F/O )
  );
  X_BUF \key2<24>1181_F/LUT4_L_BUF  (
    .I(\key2<24>1181_F/O ),
    .O(N5706)
  );
  defparam \key2<24>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<24>1181_F  (
    .ADR0(roundsel[2]),
    .ADR1(CHOICE423),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out24 ),
    .O(\key2<24>1181_F/O )
  );
  X_BUF \key2<48>961_F/LUT4_L_BUF  (
    .I(\key2<48>961_F/O ),
    .O(N5708)
  );
  defparam \key2<48>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<48>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out6 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out21 ),
    .O(\key2<48>961_F/O )
  );
  X_BUF \key2<36>1181_F/LUT4_L_BUF  (
    .I(\key2<36>1181_F/O ),
    .O(N5710)
  );
  defparam \key2<36>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<36>1181_F  (
    .ADR0(roundsel[2]),
    .ADR1(CHOICE391),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out9 ),
    .O(\key2<36>1181_F/O )
  );
  X_BUF \key2<23>1181_F/LUT4_L_BUF  (
    .I(\key2<23>1181_F/O ),
    .O(N5712)
  );
  defparam \key2<23>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<23>1181_F  (
    .ADR0(roundsel_2_7),
    .ADR1(CHOICE900),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .O(\key2<23>1181_F/O )
  );
  X_BUF \key2<48>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<48>110_SW01_F/O ),
    .O(N5714)
  );
  defparam \key2<48>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<48>110_SW01_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out55 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out31 ),
    .O(\key2<48>110_SW01_F/O )
  );
  X_BUF \c1/Mxor_X_Result<0>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_X_Result<0>11_F/O ),
    .O(N5716)
  );
  defparam \c1/Mxor_X_Result<0>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_X_Result<0>11_F  (
    .ADR0(roundsel[3]),
    .ADR1(data1[1]),
    .ADR2(CHOICE1093),
    .ADR3(\MUX_BLOCK_roundsel<2>_mmx_out33 ),
    .O(\c1/Mxor_X_Result<0>11_F/O )
  );
  X_BUF \key2<1>271_F/LUT4_L_BUF  (
    .I(\key2<1>271_F/O ),
    .O(N5718)
  );
  defparam \key2<1>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<1>271_F  (
    .ADR0(roundsel_3_16),
    .ADR1(\key1[20] ),
    .ADR2(roundsel[2]),
    .ADR3(\key1[53] ),
    .O(\key2<1>271_F/O )
  );
  X_BUF \key2<44>961_F/LUT4_L_BUF  (
    .I(\key2<44>961_F/O ),
    .O(N5720)
  );
  defparam \key2<44>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<44>961_F  (
    .ADR0(roundsel_3_5),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out92 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out55 ),
    .O(\key2<44>961_F/O )
  );
  X_BUF \key2<18>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<18>110_SW01_F/O ),
    .O(N5722)
  );
  defparam \key2<18>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<18>110_SW01_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out26 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out24 ),
    .O(\key2<18>110_SW01_F/O )
  );
  X_BUF \key2<36>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<36>133_SW01_F/O ),
    .O(N5724)
  );
  defparam \key2<36>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<36>133_SW01_F  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out13 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out10 ),
    .O(\key2<36>133_SW01_F/O )
  );
  X_BUF \key2<16>271_F/LUT4_L_BUF  (
    .I(\key2<16>271_F/O ),
    .O(N5726)
  );
  defparam \key2<16>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<16>271_F  (
    .ADR0(roundsel_3_8),
    .ADR1(\key1[11] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[12] ),
    .O(\key2<16>271_F/O )
  );
  X_BUF \c1/Mxor_X_Result<25>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_X_Result<25>11_F/O ),
    .O(N5728)
  );
  defparam \c1/Mxor_X_Result<25>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_X_Result<25>11_F  (
    .ADR0(roundsel_3_16),
    .ADR1(data1[16]),
    .ADR2(CHOICE1652),
    .ADR3(\MUX_BLOCK_roundsel<2>_mmx_out7 ),
    .O(\c1/Mxor_X_Result<25>11_F/O )
  );
  X_BUF \key2<14>1181_F/LUT4_L_BUF  (
    .I(\key2<14>1181_F/O ),
    .O(N5730)
  );
  defparam \key2<14>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<14>1181_F  (
    .ADR0(roundsel_3_10),
    .ADR1(CHOICE571),
    .ADR2(roundsel_4_8),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out44 ),
    .O(\key2<14>1181_F/O )
  );
  X_BUF \key2<12>761_F/LUT4_L_BUF  (
    .I(\key2<12>761_F/O ),
    .O(N5732)
  );
  defparam \key2<12>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<12>761_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out70 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .O(\key2<12>761_F/O )
  );
  X_BUF \key2<8>61_F/LUT3_L_BUF  (
    .I(\key2<8>61_F/O ),
    .O(N5734)
  );
  defparam \key2<8>61_F .INIT = 8'hE4;
  X_LUT3 \key2<8>61_F  (
    .ADR0(roundsel_11),
    .ADR1(\key1[50] ),
    .ADR2(\key1[58] ),
    .O(\key2<8>61_F/O )
  );
  X_BUF \key2<13>961_F/LUT4_L_BUF  (
    .I(\key2<13>961_F/O ),
    .O(N5736)
  );
  defparam \key2<13>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<13>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out68 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .O(\key2<13>961_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<2>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<2>11_F/O ),
    .O(N5738)
  );
  defparam \c1/Mxor_OUTR_Result<2>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<2>11_F  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[35]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_88 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_90 ),
    .O(\c1/Mxor_OUTR_Result<2>11_F/O )
  );
  X_BUF \key2<9>471_F/LUT4_L_BUF  (
    .I(\key2<9>471_F/O ),
    .O(N5740)
  );
  defparam \key2<9>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<9>471_F  (
    .ADR0(roundsel_3_2),
    .ADR1(\key1[51] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[52] ),
    .O(\key2<9>471_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<1>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<1>11_F/O ),
    .O(N5742)
  );
  defparam \c1/Mxor_OUTR_Result<1>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<1>11_F  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[34]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_108 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_110 ),
    .O(\c1/Mxor_OUTR_Result<1>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<9>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<9>11_F/O ),
    .O(N5744)
  );
  defparam \c1/Mxor_OUTR_Result<9>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<9>11_F  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[42]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_104 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_106 ),
    .O(\c1/Mxor_OUTR_Result<9>11_F/O )
  );
  X_BUF \key2<38>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<38>110_SW01_F/O ),
    .O(N5746)
  );
  defparam \key2<38>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<38>110_SW01_F  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out94 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out80 ),
    .O(\key2<38>110_SW01_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<15>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<15>11_F/O ),
    .O(N5748)
  );
  defparam \c1/Mxor_OUTR_Result<15>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<15>11_F  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[48]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_100 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_102 ),
    .O(\c1/Mxor_OUTR_Result<15>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<8>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<8>11_F/O ),
    .O(N5750)
  );
  defparam \c1/Mxor_OUTR_Result<8>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<8>11_F  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[41]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_80 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_82 ),
    .O(\c1/Mxor_OUTR_Result<8>11_F/O )
  );
  X_BUF \key2<41>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<41>110_SW01_F/O ),
    .O(N5752)
  );
  defparam \key2<41>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<41>110_SW01_F  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out86 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out84 ),
    .O(\key2<41>110_SW01_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<26>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<26>11_F/O ),
    .O(N5754)
  );
  defparam \c1/Mxor_OUTR_Result<26>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<26>11_F  (
    .ADR0(\c1/X[18] ),
    .ADR1(data1[59]),
    .ADR2(\c1/u2/Mrom_dout_inst_lut4_92 ),
    .ADR3(\c1/u2/Mrom_dout_inst_lut4_94 ),
    .O(\c1/Mxor_OUTR_Result<26>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<29>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<29>11_F/O ),
    .O(N5756)
  );
  defparam \c1/Mxor_OUTR_Result<29>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<29>11_F  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[62]),
    .ADR2(\c1/u4/Mrom_dout_inst_lut4_60 ),
    .ADR3(\c1/u4/Mrom_dout_inst_lut4_62 ),
    .O(\c1/Mxor_OUTR_Result<29>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<22>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<22>11_F/O ),
    .O(N5758)
  );
  defparam \c1/Mxor_OUTR_Result<22>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<22>11_F  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[55]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_72 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_74 ),
    .O(\c1/Mxor_OUTR_Result<22>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<12>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<12>11_F/O ),
    .O(N5762)
  );
  defparam \c1/Mxor_OUTR_Result<12>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<12>11_F  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[45]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_65 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_67 ),
    .O(\c1/Mxor_OUTR_Result<12>11_F/O )
  );
  X_BUF \key2<12>90_SW0_F/LUT3_L_BUF  (
    .I(\key2<12>90_SW0_F/O ),
    .O(N5764)
  );
  defparam \key2<12>90_SW0_F .INIT = 8'h27;
  X_LUT3 \key2<12>90_SW0_F  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out37 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out49 ),
    .O(\key2<12>90_SW0_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<6>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<6>11_F/O ),
    .O(N5766)
  );
  defparam \c1/Mxor_OUTR_Result<6>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<6>11_F  (
    .ADR0(\c1/X[24] ),
    .ADR1(data1[39]),
    .ADR2(\c1/u3/Mrom_dout_inst_lut4_64 ),
    .ADR3(\c1/u3/Mrom_dout_inst_lut4_66 ),
    .O(\c1/Mxor_OUTR_Result<6>11_F/O )
  );
  X_BUF \key2<46>471_F/LUT4_L_BUF  (
    .I(\key2<46>471_F/O ),
    .O(N5768)
  );
  defparam \key2<46>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<46>471_F  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[13] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[48] ),
    .O(\key2<46>471_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<27>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<27>11_F/O ),
    .O(N5770)
  );
  defparam \c1/Mxor_OUTR_Result<27>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<27>11_F  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[60]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_0 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_2 ),
    .O(\c1/Mxor_OUTR_Result<27>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<11>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<11>11_F/O ),
    .O(N5772)
  );
  defparam \c1/Mxor_OUTR_Result<11>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<11>11_F  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[44]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_12 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_14 ),
    .O(\c1/Mxor_OUTR_Result<11>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<23>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<23>11_F/O ),
    .O(N5774)
  );
  defparam \c1/Mxor_OUTR_Result<23>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<23>11_F  (
    .ADR0(\c1/X[6] ),
    .ADR1(data1[56]),
    .ADR2(\c1/u0/Mrom_dout_inst_lut4_96 ),
    .ADR3(\c1/u0/Mrom_dout_inst_lut4_98 ),
    .O(\c1/Mxor_OUTR_Result<23>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<10>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<10>11_F/O ),
    .O(N5776)
  );
  defparam \c1/Mxor_OUTR_Result<10>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<10>11_F  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[43]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_24 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_26 ),
    .O(\c1/Mxor_OUTR_Result<10>11_F/O )
  );
  X_BUF \key2<8>271_F/LUT4_L_BUF  (
    .I(\key2<8>271_F/O ),
    .O(N5778)
  );
  defparam \key2<8>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<8>271_F  (
    .ADR0(roundsel_3_8),
    .ADR1(\key1[36] ),
    .ADR2(roundsel_23),
    .ADR3(\key1[2] ),
    .O(\key2<8>271_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<5>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<5>11_F/O ),
    .O(N5780)
  );
  defparam \c1/Mxor_OUTR_Result<5>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<5>11_F  (
    .ADR0(\c1/X[48] ),
    .ADR1(data1[38]),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_4 ),
    .ADR3(\c1/u7/Mrom_dout_inst_lut4_6 ),
    .O(\c1/Mxor_OUTR_Result<5>11_F/O )
  );
  X_BUF \key2<40>761_F/LUT4_L_BUF  (
    .I(\key2<40>761_F/O ),
    .O(N5782)
  );
  defparam \key2<40>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<40>761_F  (
    .ADR0(roundsel_4_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out82 ),
    .ADR2(roundsel_3_13),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out87 ),
    .O(\key2<40>761_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<18>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<18>11_F/O ),
    .O(N5784)
  );
  defparam \c1/Mxor_OUTR_Result<18>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<18>11_F  (
    .ADR0(\c1/X[30] ),
    .ADR1(data1[51]),
    .ADR2(\c1/u4/Mrom_dout_inst_lut4_52 ),
    .ADR3(\c1/u4/Mrom_dout_inst_lut4_54 ),
    .O(\c1/Mxor_OUTR_Result<18>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<0>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<0>11_F/O ),
    .O(N5786)
  );
  defparam \c1/Mxor_OUTR_Result<0>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<0>11_F  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[33]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_16 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_18 ),
    .O(\c1/Mxor_OUTR_Result<0>11_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<17>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<17>11_F/O ),
    .O(N5788)
  );
  defparam \c1/Mxor_OUTR_Result<17>11_F .INIT = 16'h6A59;
  X_LUT4 \c1/Mxor_OUTR_Result<17>11_F  (
    .ADR0(data1[50]),
    .ADR1(\c1/X[48] ),
    .ADR2(\c1/u7/Mrom_dout_inst_lut4_10 ),
    .ADR3(N5490),
    .O(\c1/Mxor_OUTR_Result<17>11_F/O )
  );
  X_BUF \key2<2>961_F/LUT4_L_BUF  (
    .I(\key2<2>961_F/O ),
    .O(N5790)
  );
  defparam \key2<2>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<2>961_F  (
    .ADR0(roundsel_3_5),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out42 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out67 ),
    .O(\key2<2>961_F/O )
  );
  X_BUF \key2<26>271_F/LUT4_L_BUF  (
    .I(\key2<26>271_F/O ),
    .O(N5792)
  );
  defparam \key2<26>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<26>271_F  (
    .ADR0(roundsel_3_7),
    .ADR1(\key1[29] ),
    .ADR2(roundsel_22),
    .ADR3(\key1[64] ),
    .O(\key2<26>271_F/O )
  );
  X_BUF \key2<29>1181_F/LUT4_L_BUF  (
    .I(\key2<29>1181_F/O ),
    .O(N5794)
  );
  defparam \key2<29>1181_F .INIT = 16'h0E04;
  X_LUT4 \key2<29>1181_F  (
    .ADR0(roundsel_4_3),
    .ADR1(CHOICE1545),
    .ADR2(roundsel_3_14),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out21 ),
    .O(\key2<29>1181_F/O )
  );
  X_BUF \key2<15>1191_F/LUT4_L_BUF  (
    .I(\key2<15>1191_F/O ),
    .O(N5796)
  );
  defparam \key2<15>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<15>1191_F  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out53 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out25 ),
    .O(\key2<15>1191_F/O )
  );
  X_BUF \key2<20>961_F/LUT4_L_BUF  (
    .I(\key2<20>961_F/O ),
    .O(N5798)
  );
  defparam \key2<20>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<20>961_F  (
    .ADR0(roundsel_3_13),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out46 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out48 ),
    .O(\key2<20>961_F/O )
  );
  X_BUF \key2<37>271_F/LUT4_L_BUF  (
    .I(\key2<37>271_F/O ),
    .O(N5800)
  );
  defparam \key2<37>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<37>271_F  (
    .ADR0(roundsel_33),
    .ADR1(\key1[5] ),
    .ADR2(roundsel_2_13),
    .ADR3(\key1[40] ),
    .O(\key2<37>271_F/O )
  );
  X_BUF \key2<11>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<11>110_SW01_F/O ),
    .O(N5802)
  );
  defparam \key2<11>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<11>110_SW01_F  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out60 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out29 ),
    .O(\key2<11>110_SW01_F/O )
  );
  X_BUF \key2<25>271_F/LUT4_L_BUF  (
    .I(\key2<25>271_F/O ),
    .O(N5804)
  );
  defparam \key2<25>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<25>271_F  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[6] ),
    .ADR2(roundsel_2_4),
    .ADR3(\key1[5] ),
    .O(\key2<25>271_F/O )
  );
  X_BUF \key2<11>961_F/LUT4_L_BUF  (
    .I(\key2<11>961_F/O ),
    .O(N5806)
  );
  defparam \key2<11>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<11>961_F  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out63 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out65 ),
    .O(\key2<11>961_F/O )
  );
  X_BUF \key2<39>90_SW01_F/LUT3_L_BUF  (
    .I(\key2<39>90_SW01_F/O ),
    .O(N5808)
  );
  defparam \key2<39>90_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<39>90_SW01_F  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out31 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out77 ),
    .O(\key2<39>90_SW01_F/O )
  );
  X_BUF \key2<23>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<23>133_SW01_F/O ),
    .O(N5810)
  );
  defparam \key2<23>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<23>133_SW01_F  (
    .ADR0(roundsel_2_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out33 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out32 ),
    .O(\key2<23>133_SW01_F/O )
  );
  X_BUF \key2<30>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<30>133_SW01_F/O ),
    .O(N5812)
  );
  defparam \key2<30>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<30>133_SW01_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out91 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out20 ),
    .O(\key2<30>133_SW01_F/O )
  );
  X_BUF \key2<46>1191_F/LUT4_L_BUF  (
    .I(\key2<46>1191_F/O ),
    .O(N5814)
  );
  defparam \key2<46>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<46>1191_F  (
    .ADR0(roundsel_3_13),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out83 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out85 ),
    .O(\key2<46>1191_F/O )
  );
  X_BUF \key2<13>271_F/LUT4_L_BUF  (
    .I(\key2<13>271_F/O ),
    .O(N5816)
  );
  defparam \key2<13>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<13>271_F  (
    .ADR0(roundsel_33),
    .ADR1(\key1[50] ),
    .ADR2(roundsel_2_10),
    .ADR3(\key1[51] ),
    .O(\key2<13>271_F/O )
  );
  X_BUF \key2<42>961_F/LUT4_L_BUF  (
    .I(\key2<42>961_F/O ),
    .O(N5818)
  );
  defparam \key2<42>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<42>961_F  (
    .ADR0(roundsel[3]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out4 ),
    .ADR2(roundsel[4]),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out91 ),
    .O(\key2<42>961_F/O )
  );
  X_BUF \key2<10>961_F/LUT4_L_BUF  (
    .I(\key2<10>961_F/O ),
    .O(N5820)
  );
  defparam \key2<10>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<10>961_F  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out30 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out34 ),
    .O(\key2<10>961_F/O )
  );
  X_BUF \key2<15>471_F/LUT4_L_BUF  (
    .I(\key2<15>471_F/O ),
    .O(N5822)
  );
  defparam \key2<15>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<15>471_F  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[26] ),
    .ADR2(roundsel_3_1),
    .ADR3(\key1[58] ),
    .O(\key2<15>471_F/O )
  );
  X_BUF \key2<9>1191_F/LUT4_L_BUF  (
    .I(\key2<9>1191_F/O ),
    .O(N5824)
  );
  defparam \key2<9>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<9>1191_F  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out58 ),
    .ADR2(roundsel_43),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out29 ),
    .O(\key2<9>1191_F/O )
  );
  X_BUF \key2<27>471_F/LUT4_L_BUF  (
    .I(\key2<27>471_F/O ),
    .O(N5826)
  );
  defparam \key2<27>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<27>471_F  (
    .ADR0(roundsel_3_1),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_2_1),
    .ADR3(\key1[55] ),
    .O(\key2<27>471_F/O )
  );
  X_BUF \c1/Mxor_X_Result<31>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_X_Result<31>11_F/O ),
    .O(N5828)
  );
  defparam \c1/Mxor_X_Result<31>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_X_Result<31>11_F  (
    .ADR0(roundsel_3_14),
    .ADR1(data1[12]),
    .ADR2(CHOICE1676),
    .ADR3(\MUX_BLOCK_roundsel<2>_mmx_out11 ),
    .O(\c1/Mxor_X_Result<31>11_F/O )
  );
  X_BUF \key2<24>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<24>133_SW01_F/O ),
    .O(N5830)
  );
  defparam \key2<24>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<24>133_SW01_F  (
    .ADR0(roundsel[2]),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out28 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .O(\key2<24>133_SW01_F/O )
  );
  X_BUF \key2<27>1411_F/LUT4_L_BUF  (
    .I(\key2<27>1411_F/O ),
    .O(N5832)
  );
  defparam \key2<27>1411_F .INIT = 16'h0E04;
  X_LUT4 \key2<27>1411_F  (
    .ADR0(roundsel_3_5),
    .ADR1(CHOICE1332),
    .ADR2(roundsel_4_7),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out90 ),
    .O(\key2<27>1411_F/O )
  );
  X_BUF \key2<10>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<10>110_SW01_F/O ),
    .O(N5834)
  );
  defparam \key2<10>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<10>110_SW01_F  (
    .ADR0(roundsel_3_3),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out50 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out41 ),
    .O(\key2<10>110_SW01_F/O )
  );
  X_BUF \key2<2>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<2>110_SW01_F/O ),
    .O(N5836)
  );
  defparam \key2<2>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<2>110_SW01_F  (
    .ADR0(roundsel_3_11),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out45 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out60 ),
    .O(\key2<2>110_SW01_F/O )
  );
  X_BUF \key2<5>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<5>110_SW01_F/O ),
    .O(N5838)
  );
  defparam \key2<5>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<5>110_SW01_F  (
    .ADR0(roundsel_2_7),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out72 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out65 ),
    .O(\key2<5>110_SW01_F/O )
  );
  X_BUF \key2<7>761_F/LUT4_L_BUF  (
    .I(\key2<7>761_F/O ),
    .O(N5840)
  );
  defparam \key2<7>761_F .INIT = 16'h0E04;
  X_LUT4 \key2<7>761_F  (
    .ADR0(roundsel_33),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out56 ),
    .ADR2(roundsel_4_5),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out72 ),
    .O(\key2<7>761_F/O )
  );
  X_BUF \key2<33>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<33>110_SW01_F/O ),
    .O(N5842)
  );
  defparam \key2<33>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<33>110_SW01_F  (
    .ADR0(roundsel_3_2),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out9 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out85 ),
    .O(\key2<33>110_SW01_F/O )
  );
  X_BUF \key2<45>1191_F/LUT4_L_BUF  (
    .I(\key2<45>1191_F/O ),
    .O(N5844)
  );
  defparam \key2<45>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<45>1191_F  (
    .ADR0(roundsel_23),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out89 ),
    .ADR2(roundsel_3_13),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out90 ),
    .O(\key2<45>1191_F/O )
  );
  X_BUF \key2<5>961_F/LUT4_L_BUF  (
    .I(\key2<5>961_F/O ),
    .O(N5846)
  );
  defparam \key2<5>961_F .INIT = 16'h0E04;
  X_LUT4 \key2<5>961_F  (
    .ADR0(roundsel_2_6),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out71 ),
    .ADR2(roundsel_4_6),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out38 ),
    .O(\key2<5>961_F/O )
  );
  X_BUF \key2<14>133_SW01_F/LUT3_L_BUF  (
    .I(\key2<14>133_SW01_F/O ),
    .O(N5848)
  );
  defparam \key2<14>133_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<14>133_SW01_F  (
    .ADR0(roundsel_3_12),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out27 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out61 ),
    .O(\key2<14>133_SW01_F/O )
  );
  X_BUF \key2<43>271_F/LUT4_L_BUF  (
    .I(\key2<43>271_F/O ),
    .O(N5850)
  );
  defparam \key2<43>271_F .INIT = 16'h0E04;
  X_LUT4 \key2<43>271_F  (
    .ADR0(roundsel_33),
    .ADR1(\key1[30] ),
    .ADR2(roundsel_2_10),
    .ADR3(\key1[29] ),
    .O(\key2<43>271_F/O )
  );
  X_BUF \c1/Mxor_X_Result<15>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_X_Result<15>11_F/O ),
    .O(N5852)
  );
  defparam \c1/Mxor_X_Result<15>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_X_Result<15>11_F  (
    .ADR0(roundsel_3_16),
    .ADR1(data1[22]),
    .ADR2(CHOICE510),
    .ADR3(\MUX_BLOCK_roundsel<2>_mmx_out27 ),
    .O(\c1/Mxor_X_Result<15>11_F/O )
  );
  X_BUF \key2<28>471_F/LUT4_L_BUF  (
    .I(\key2<28>471_F/O ),
    .O(N5854)
  );
  defparam \key2<28>471_F .INIT = 16'h0E04;
  X_LUT4 \key2<28>471_F  (
    .ADR0(roundsel_2_1),
    .ADR1(\key1[56] ),
    .ADR2(roundsel_4_1),
    .ADR3(\key1[23] ),
    .O(\key2<28>471_F/O )
  );
  X_BUF \key2<17>1191_F/LUT4_L_BUF  (
    .I(\key2<17>1191_F/O ),
    .O(N5856)
  );
  defparam \key2<17>1191_F .INIT = 16'h0E04;
  X_LUT4 \key2<17>1191_F  (
    .ADR0(roundsel_2_8),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out59 ),
    .ADR2(roundsel_4_9),
    .ADR3(\MUX_BLOCK_roundsel<1>_mmx_out60 ),
    .O(\key2<17>1191_F/O )
  );
  X_BUF \key2<20>110_SW01_F/LUT3_L_BUF  (
    .I(\key2<20>110_SW01_F/O ),
    .O(N5858)
  );
  defparam \key2<20>110_SW01_F .INIT = 8'h27;
  X_LUT3 \key2<20>110_SW01_F  (
    .ADR0(roundsel_3_15),
    .ADR1(\MUX_BLOCK_roundsel<1>_mmx_out52 ),
    .ADR2(\MUX_BLOCK_roundsel<1>_mmx_out50 ),
    .O(\key2<20>110_SW01_F/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_291_F/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_291_F/O ),
    .O(N5860)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_291_F .INIT = 16'h9D61;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_291_F  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[27] ),
    .ADR2(\c1/X[28] ),
    .ADR3(\c1/X[29] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_291_F/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_281_F/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_281_F/O ),
    .O(N5862)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_281_F .INIT = 16'h693C;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_281_F  (
    .ADR0(\c1/X[29] ),
    .ADR1(\c1/X[26] ),
    .ADR2(\c1/X[28] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_281_F/O )
  );
  X_BUF \roundsel<2>_mmx_out331_F/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out331_F/O ),
    .O(N5864)
  );
  defparam \roundsel<2>_mmx_out331_F .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out331_F  (
    .ADR0(roundsel_1_3),
    .ADR1(\key1[27] ),
    .ADR2(\key1[43] ),
    .O(\roundsel<2>_mmx_out331_F/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_251_F/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_251_F/O ),
    .O(N5866)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_251_F .INIT = 16'h26BC;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_251_F  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[27] ),
    .ADR2(\c1/X[29] ),
    .ADR3(\c1/X[28] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_251_F/O )
  );
  X_BUF \c1/u4/Mrom_dout_inst_mux_f5_241_F/LUT4_L_BUF  (
    .I(\c1/u4/Mrom_dout_inst_mux_f5_241_F/O ),
    .O(N5868)
  );
  defparam \c1/u4/Mrom_dout_inst_mux_f5_241_F .INIT = 16'hB664;
  X_LUT4 \c1/u4/Mrom_dout_inst_mux_f5_241_F  (
    .ADR0(\c1/X[26] ),
    .ADR1(\c1/X[28] ),
    .ADR2(\c1/X[29] ),
    .ADR3(\c1/X[27] ),
    .O(\c1/u4/Mrom_dout_inst_mux_f5_241_F/O )
  );
  X_BUF \c1/u6/Mrom_dout_inst_mux_f5_111_F/LUT4_L_BUF  (
    .I(\c1/u6/Mrom_dout_inst_mux_f5_111_F/O ),
    .O(N5870)
  );
  defparam \c1/u6/Mrom_dout_inst_mux_f5_111_F .INIT = 16'hA674;
  X_LUT4 \c1/u6/Mrom_dout_inst_mux_f5_111_F  (
    .ADR0(\c1/X[40] ),
    .ADR1(\c1/X[41] ),
    .ADR2(\c1/X[39] ),
    .ADR3(\c1/X[38] ),
    .O(\c1/u6/Mrom_dout_inst_mux_f5_111_F/O )
  );
  X_BUF \c1/u6/Mrom_dout_inst_mux_f5_101_F/LUT4_L_BUF  (
    .I(\c1/u6/Mrom_dout_inst_mux_f5_101_F/O ),
    .O(N5872)
  );
  defparam \c1/u6/Mrom_dout_inst_mux_f5_101_F .INIT = 16'h6396;
  X_LUT4 \c1/u6/Mrom_dout_inst_mux_f5_101_F  (
    .ADR0(\c1/X[39] ),
    .ADR1(\c1/X[40] ),
    .ADR2(\c1/X[41] ),
    .ADR3(\c1/X[38] ),
    .O(\c1/u6/Mrom_dout_inst_mux_f5_101_F/O )
  );
  X_BUF \c1/Mxor_OUTR_Result<25>11_F/LUT4_L_BUF  (
    .I(\c1/Mxor_OUTR_Result<25>11_F/O ),
    .O(N5874)
  );
  defparam \c1/Mxor_OUTR_Result<25>11_F .INIT = 16'h369C;
  X_LUT4 \c1/Mxor_OUTR_Result<25>11_F  (
    .ADR0(\c1/X[42] ),
    .ADR1(data1[58]),
    .ADR2(\c1/u6/Mrom_dout_inst_lut4_26 ),
    .ADR3(\c1/u6/Mrom_dout_inst_lut4_30 ),
    .O(\c1/Mxor_OUTR_Result<25>11_F/O )
  );
  X_BUF \roundsel<2>_mmx_out241_F/LUT3_L_BUF  (
    .I(\roundsel<2>_mmx_out241_F/O ),
    .O(N5876)
  );
  defparam \roundsel<2>_mmx_out241_F .INIT = 8'hE4;
  X_LUT3 \roundsel<2>_mmx_out241_F  (
    .ADR0(roundsel_12),
    .ADR1(\key1[43] ),
    .ADR2(\key1[59] ),
    .O(\roundsel<2>_mmx_out241_F/O )
  );
  X_BUF \key2<31>15_F/LUT4_L_BUF  (
    .I(\key2<31>15_F/O ),
    .O(N5878)
  );
  defparam \key2<31>15_F .INIT = 16'h0E04;
  X_LUT4 \key2<31>15_F  (
    .ADR0(roundsel_1_20),
    .ADR1(\key1[54] ),
    .ADR2(roundsel_3_16),
    .ADR3(\key1[5] ),
    .O(\key2<31>15_F/O )
  );
  X_BUF \key2<26>12_F/LUT4_L_BUF  (
    .I(\key2<26>12_F/O ),
    .O(N5880)
  );
  defparam \key2<26>12_F .INIT = 16'hA280;
  X_LUT4 \key2<26>12_F  (
    .ADR0(roundsel_2_6),
    .ADR1(roundsel_1_17),
    .ADR2(\key1[48] ),
    .ADR3(\key1[32] ),
    .O(\key2<26>12_F/O )
  );
  X_BUF \key2<8>12_F/LUT4_L_BUF  (
    .I(\key2<8>12_F/O ),
    .O(N5882)
  );
  defparam \key2<8>12_F .INIT = 16'hA280;
  X_LUT4 \key2<8>12_F  (
    .ADR0(roundsel_2_8),
    .ADR1(roundsel_1_4),
    .ADR2(\key1[53] ),
    .ADR3(\key1[37] ),
    .O(\key2<8>12_F/O )
  );
  X_BUF \key2<37>12_SW0_F/LUT3_L_BUF  (
    .I(\key2<37>12_SW0_F/O ),
    .O(N5884)
  );
  defparam \key2<37>12_SW0_F .INIT = 8'hE4;
  X_LUT3 \key2<37>12_SW0_F  (
    .ADR0(roundsel_11),
    .ADR1(\key1[8] ),
    .ADR2(\key1[24] ),
    .O(\key2<37>12_SW0_F/O )
  );
  X_BUF \key2<43>12_SW0_F/LUT3_L_BUF  (
    .I(\key2<43>12_SW0_F/O ),
    .O(N5886)
  );
  defparam \key2<43>12_SW0_F .INIT = 8'hE4;
  X_LUT3 \key2<43>12_SW0_F  (
    .ADR0(roundsel_11),
    .ADR1(\key1[62] ),
    .ADR2(\key1[13] ),
    .O(\key2<43>12_SW0_F/O )
  );
  X_BUF \key2<13>12_SW0_F/LUT3_L_BUF  (
    .I(\key2<13>12_SW0_F/O ),
    .O(N5888)
  );
  defparam \key2<13>12_SW0_F .INIT = 8'hE4;
  X_LUT3 \key2<13>12_SW0_F  (
    .ADR0(roundsel_1_3),
    .ADR1(\key1[19] ),
    .ADR2(\key1[35] ),
    .O(\key2<13>12_SW0_F/O )
  );
  X_BUF \key2<7>15_F/LUT4_L_BUF  (
    .I(\key2<7>15_F/O ),
    .O(N5890)
  );
  defparam \key2<7>15_F .INIT = 16'h0E04;
  X_LUT4 \key2<7>15_F  (
    .ADR0(roundsel_12),
    .ADR1(\key1[27] ),
    .ADR2(roundsel_3_6),
    .ADR3(\key1[43] ),
    .O(\key2<7>15_F/O )
  );
  X_BUF \key2<26>61_F/LUT3_L_BUF  (
    .I(\key2<26>61_F/O ),
    .O(N5892)
  );
  defparam \key2<26>61_F .INIT = 8'hE4;
  X_LUT3 \key2<26>61_F  (
    .ADR0(roundsel_1_11),
    .ADR1(\key1[47] ),
    .ADR2(\key1[55] ),
    .O(\key2<26>61_F/O )
  );
  X_BUF \key2<31>12_F/LUT4_L_BUF  (
    .I(\key2<31>12_F/O ),
    .O(N5894)
  );
  defparam \key2<31>12_F .INIT = 16'hA280;
  X_LUT4 \key2<31>12_F  (
    .ADR0(roundsel_3_6),
    .ADR1(roundsel_1_2),
    .ADR2(\key1[40] ),
    .ADR3(\key1[24] ),
    .O(\key2<31>12_F/O )
  );
  X_CKBUF \clk_BUFGP/BUFG  (
    .I(\clk_BUFGP/IBUFG ),
    .O(clk_BUFGP)
  );
  X_CKBUF \clk_BUFGP/IBUFG_252  (
    .I(clk),
    .O(\clk_BUFGP/IBUFG )
  );
  X_TRI \dataout_1_OBUF.GTS.TRI_253  (
    .I(\dataout_1_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_1_OBUF.GTS.TRI/CTL ),
    .O(dataout[1])
  );
  X_TRI \dataout_23_OBUF.GTS.TRI_254  (
    .I(\dataout_23_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_23_OBUF.GTS.TRI/CTL ),
    .O(dataout[23])
  );
  X_TRI \dataout_4_OBUF.GTS.TRI_255  (
    .I(\dataout_4_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_4_OBUF.GTS.TRI/CTL ),
    .O(dataout[4])
  );
  X_TRI \dataout_48_OBUF.GTS.TRI_256  (
    .I(\dataout_48_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_48_OBUF.GTS.TRI/CTL ),
    .O(dataout[48])
  );
  X_TRI \dataout_43_OBUF.GTS.TRI_257  (
    .I(\dataout_43_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_43_OBUF.GTS.TRI/CTL ),
    .O(dataout[43])
  );
  X_TRI \dataout_25_OBUF.GTS.TRI_258  (
    .I(\dataout_25_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_25_OBUF.GTS.TRI/CTL ),
    .O(dataout[25])
  );
  X_TRI \dataout_49_OBUF.GTS.TRI_259  (
    .I(\dataout_49_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_49_OBUF.GTS.TRI/CTL ),
    .O(dataout[49])
  );
  X_TRI \dataout_31_OBUF.GTS.TRI_260  (
    .I(\dataout_31_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_31_OBUF.GTS.TRI/CTL ),
    .O(dataout[31])
  );
  X_TRI \dataout_24_OBUF.GTS.TRI_261  (
    .I(\dataout_24_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_24_OBUF.GTS.TRI/CTL ),
    .O(dataout[24])
  );
  X_TRI \dataout_35_OBUF.GTS.TRI_262  (
    .I(\dataout_35_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_35_OBUF.GTS.TRI/CTL ),
    .O(dataout[35])
  );
  X_TRI \dataout_33_OBUF.GTS.TRI_263  (
    .I(\dataout_33_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_33_OBUF.GTS.TRI/CTL ),
    .O(dataout[33])
  );
  X_TRI \dataout_46_OBUF.GTS.TRI_264  (
    .I(\dataout_46_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_46_OBUF.GTS.TRI/CTL ),
    .O(dataout[46])
  );
  X_TRI \dataout_26_OBUF.GTS.TRI_265  (
    .I(\dataout_26_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_26_OBUF.GTS.TRI/CTL ),
    .O(dataout[26])
  );
  X_TRI \dataout_17_OBUF.GTS.TRI_266  (
    .I(\dataout_17_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_17_OBUF.GTS.TRI/CTL ),
    .O(dataout[17])
  );
  X_TRI \dataout_45_OBUF.GTS.TRI_267  (
    .I(\dataout_45_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_45_OBUF.GTS.TRI/CTL ),
    .O(dataout[45])
  );
  X_TRI \dataout_40_OBUF.GTS.TRI_268  (
    .I(\dataout_40_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_40_OBUF.GTS.TRI/CTL ),
    .O(dataout[40])
  );
  X_TRI \dataout_42_OBUF.GTS.TRI_269  (
    .I(\dataout_42_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_42_OBUF.GTS.TRI/CTL ),
    .O(dataout[42])
  );
  X_TRI \dataout_6_OBUF.GTS.TRI_270  (
    .I(\dataout_6_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_6_OBUF.GTS.TRI/CTL ),
    .O(dataout[6])
  );
  X_TRI \dataout_3_OBUF.GTS.TRI_271  (
    .I(\dataout_3_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_3_OBUF.GTS.TRI/CTL ),
    .O(dataout[3])
  );
  X_TRI \dataout_51_OBUF.GTS.TRI_272  (
    .I(\dataout_51_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_51_OBUF.GTS.TRI/CTL ),
    .O(dataout[51])
  );
  X_TRI \dataout_28_OBUF.GTS.TRI_273  (
    .I(\dataout_28_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_28_OBUF.GTS.TRI/CTL ),
    .O(dataout[28])
  );
  X_TRI \dataout_5_OBUF.GTS.TRI_274  (
    .I(\dataout_5_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_5_OBUF.GTS.TRI/CTL ),
    .O(dataout[5])
  );
  X_TRI \dataout_37_OBUF.GTS.TRI_275  (
    .I(\dataout_37_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_37_OBUF.GTS.TRI/CTL ),
    .O(dataout[37])
  );
  X_TRI \dataout_36_OBUF.GTS.TRI_276  (
    .I(\dataout_36_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_36_OBUF.GTS.TRI/CTL ),
    .O(dataout[36])
  );
  X_TRI \dataout_30_OBUF.GTS.TRI_277  (
    .I(\dataout_30_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_30_OBUF.GTS.TRI/CTL ),
    .O(dataout[30])
  );
  X_TRI \dataout_39_OBUF.GTS.TRI_278  (
    .I(\dataout_39_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_39_OBUF.GTS.TRI/CTL ),
    .O(dataout[39])
  );
  X_TRI \dataout_32_OBUF.GTS.TRI_279  (
    .I(\dataout_32_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_32_OBUF.GTS.TRI/CTL ),
    .O(dataout[32])
  );
  X_TRI \dataout_29_OBUF.GTS.TRI_280  (
    .I(\dataout_29_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_29_OBUF.GTS.TRI/CTL ),
    .O(dataout[29])
  );
  X_TRI \dataout_27_OBUF.GTS.TRI_281  (
    .I(\dataout_27_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_27_OBUF.GTS.TRI/CTL ),
    .O(dataout[27])
  );
  X_TRI \dataout_34_OBUF.GTS.TRI_282  (
    .I(\dataout_34_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_34_OBUF.GTS.TRI/CTL ),
    .O(dataout[34])
  );
  X_TRI \dataout_47_OBUF.GTS.TRI_283  (
    .I(\dataout_47_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_47_OBUF.GTS.TRI/CTL ),
    .O(dataout[47])
  );
  X_TRI \dataout_38_OBUF.GTS.TRI_284  (
    .I(\dataout_38_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_38_OBUF.GTS.TRI/CTL ),
    .O(dataout[38])
  );
  X_TRI \dataout_41_OBUF.GTS.TRI_285  (
    .I(\dataout_41_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_41_OBUF.GTS.TRI/CTL ),
    .O(dataout[41])
  );
  X_TRI \dataout_50_OBUF.GTS.TRI_286  (
    .I(\dataout_50_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_50_OBUF.GTS.TRI/CTL ),
    .O(dataout[50])
  );
  X_TRI \dataout_44_OBUF.GTS.TRI_287  (
    .I(\dataout_44_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_44_OBUF.GTS.TRI/CTL ),
    .O(dataout[44])
  );
  X_TRI \dataout_2_OBUF.GTS.TRI_288  (
    .I(\dataout_2_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_2_OBUF.GTS.TRI/CTL ),
    .O(dataout[2])
  );
  X_TRI \ready_OBUF.GTS.TRI_289  (
    .I(\ready_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_ready_OBUF.GTS.TRI/CTL ),
    .O(ready)
  );
  X_TRI \dataout_15_OBUF.GTS.TRI_290  (
    .I(\dataout_15_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_15_OBUF.GTS.TRI/CTL ),
    .O(dataout[15])
  );
  X_TRI \dataout_11_OBUF.GTS.TRI_291  (
    .I(\dataout_11_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_11_OBUF.GTS.TRI/CTL ),
    .O(dataout[11])
  );
  X_TRI \dataout_14_OBUF.GTS.TRI_292  (
    .I(\dataout_14_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_14_OBUF.GTS.TRI/CTL ),
    .O(dataout[14])
  );
  X_TRI \dataout_61_OBUF.GTS.TRI_293  (
    .I(\dataout_61_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_61_OBUF.GTS.TRI/CTL ),
    .O(dataout[61])
  );
  X_TRI \dataout_7_OBUF.GTS.TRI_294  (
    .I(\dataout_7_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_7_OBUF.GTS.TRI/CTL ),
    .O(dataout[7])
  );
  X_TRI \dataout_63_OBUF.GTS.TRI_295  (
    .I(\dataout_63_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_63_OBUF.GTS.TRI/CTL ),
    .O(dataout[63])
  );
  X_TRI \dataout_64_OBUF.GTS.TRI_296  (
    .I(\dataout_64_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_64_OBUF.GTS.TRI/CTL ),
    .O(dataout[64])
  );
  X_TRI \dataout_8_OBUF.GTS.TRI_297  (
    .I(\dataout_8_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_8_OBUF.GTS.TRI/CTL ),
    .O(dataout[8])
  );
  X_TRI \dataout_52_OBUF.GTS.TRI_298  (
    .I(\dataout_52_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_52_OBUF.GTS.TRI/CTL ),
    .O(dataout[52])
  );
  X_TRI \dataout_9_OBUF.GTS.TRI_299  (
    .I(\dataout_9_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_9_OBUF.GTS.TRI/CTL ),
    .O(dataout[9])
  );
  X_TRI \dataout_56_OBUF.GTS.TRI_300  (
    .I(\dataout_56_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_56_OBUF.GTS.TRI/CTL ),
    .O(dataout[56])
  );
  X_TRI \dataout_21_OBUF.GTS.TRI_301  (
    .I(\dataout_21_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_21_OBUF.GTS.TRI/CTL ),
    .O(dataout[21])
  );
  X_TRI \dataout_62_OBUF.GTS.TRI_302  (
    .I(\dataout_62_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_62_OBUF.GTS.TRI/CTL ),
    .O(dataout[62])
  );
  X_TRI \dataout_57_OBUF.GTS.TRI_303  (
    .I(\dataout_57_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_57_OBUF.GTS.TRI/CTL ),
    .O(dataout[57])
  );
  X_TRI \dataout_19_OBUF.GTS.TRI_304  (
    .I(\dataout_19_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_19_OBUF.GTS.TRI/CTL ),
    .O(dataout[19])
  );
  X_TRI \dataout_60_OBUF.GTS.TRI_305  (
    .I(\dataout_60_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_60_OBUF.GTS.TRI/CTL ),
    .O(dataout[60])
  );
  X_TRI \dataout_58_OBUF.GTS.TRI_306  (
    .I(\dataout_58_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_58_OBUF.GTS.TRI/CTL ),
    .O(dataout[58])
  );
  X_TRI \dataout_10_OBUF.GTS.TRI_307  (
    .I(\dataout_10_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_10_OBUF.GTS.TRI/CTL ),
    .O(dataout[10])
  );
  X_TRI \dataout_55_OBUF.GTS.TRI_308  (
    .I(\dataout_55_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_55_OBUF.GTS.TRI/CTL ),
    .O(dataout[55])
  );
  X_TRI \dataout_54_OBUF.GTS.TRI_309  (
    .I(\dataout_54_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_54_OBUF.GTS.TRI/CTL ),
    .O(dataout[54])
  );
  X_TRI \dataout_12_OBUF.GTS.TRI_310  (
    .I(\dataout_12_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_12_OBUF.GTS.TRI/CTL ),
    .O(dataout[12])
  );
  X_TRI \dataout_22_OBUF.GTS.TRI_311  (
    .I(\dataout_22_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_22_OBUF.GTS.TRI/CTL ),
    .O(dataout[22])
  );
  X_TRI \dataout_16_OBUF.GTS.TRI_312  (
    .I(\dataout_16_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_16_OBUF.GTS.TRI/CTL ),
    .O(dataout[16])
  );
  X_TRI \dataout_59_OBUF.GTS.TRI_313  (
    .I(\dataout_59_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_59_OBUF.GTS.TRI/CTL ),
    .O(dataout[59])
  );
  X_TRI \dataout_13_OBUF.GTS.TRI_314  (
    .I(\dataout_13_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_13_OBUF.GTS.TRI/CTL ),
    .O(dataout[13])
  );
  X_TRI \dataout_18_OBUF.GTS.TRI_315  (
    .I(\dataout_18_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_18_OBUF.GTS.TRI/CTL ),
    .O(dataout[18])
  );
  X_TRI \dataout_53_OBUF.GTS.TRI_316  (
    .I(\dataout_53_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_53_OBUF.GTS.TRI/CTL ),
    .O(dataout[53])
  );
  X_TRI \dataout_20_OBUF.GTS.TRI_317  (
    .I(\dataout_20_OBUF.GTS.TRI ),
    .CTL(\NlwInverterSignal_dataout_20_OBUF.GTS.TRI/CTL ),
    .O(dataout[20])
  );
  X_ONE NlwBlock_des_VCC (
    .O(VCC)
  );
  X_ZERO NlwBlock_des_GND (
    .O(GND)
  );
  X_INV \NlwInverterBlock_dataout_1_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_1_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_23_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_23_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_4_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_4_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_48_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_48_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_43_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_43_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_25_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_25_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_49_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_49_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_31_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_31_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_24_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_24_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_35_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_35_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_33_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_33_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_46_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_46_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_26_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_26_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_17_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_17_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_45_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_45_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_40_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_40_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_42_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_42_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_6_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_6_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_3_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_3_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_51_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_51_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_28_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_28_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_5_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_5_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_37_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_37_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_36_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_36_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_30_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_30_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_39_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_39_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_32_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_32_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_29_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_29_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_27_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_27_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_34_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_34_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_47_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_47_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_38_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_38_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_41_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_41_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_50_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_50_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_44_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_44_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_2_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_2_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_ready_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_ready_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_15_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_15_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_11_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_11_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_14_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_14_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_61_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_61_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_7_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_7_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_63_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_63_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_64_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_64_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_8_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_8_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_52_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_52_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_9_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_9_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_56_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_56_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_21_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_21_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_62_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_62_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_57_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_57_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_19_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_19_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_60_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_60_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_58_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_58_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_10_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_10_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_55_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_55_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_54_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_54_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_12_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_12_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_22_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_22_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_16_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_16_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_59_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_59_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_13_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_13_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_18_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_18_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_53_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_53_OBUF.GTS.TRI/CTL )
  );
  X_INV \NlwInverterBlock_dataout_20_OBUF.GTS.TRI/CTL  (
    .I(GTS),
    .O(\NlwInverterSignal_dataout_20_OBUF.GTS.TRI/CTL )
  );


endmodule