--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:15:19 05/03/2013
-- Design Name:   
-- Module Name:   E:/LIZI/RSA/testbench.vhd
-- Project Name:  RSA
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: RSACypher
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY testbench IS
END testbench;

ARCHITECTURE behavior OF testbench IS 

	COMPONENT ARS_rsacypher
	PORT(
		indata : IN std_logic_vector(1023 downto 0);
		inexp : IN std_logic_vector(1023 downto 0);
		inmod : IN std_logic_vector(1023 downto 0);
		clk : IN std_logic;
		ds : IN std_logic;
		reset : IN std_logic;          
		cypher : OUT std_logic_vector(1023 downto 0);
		ready : OUT std_logic
		);
	END COMPONENT;

	SIGNAL indata :  std_logic_vector(1023 downto 0);
	SIGNAL inexp :  std_logic_vector(1023 downto 0);
	SIGNAL inmod :  std_logic_vector(1023 downto 0);
	SIGNAL cypher :  std_logic_vector(1023 downto 0);
	SIGNAL clk :  std_logic;
	SIGNAL ds :  std_logic;
	SIGNAL reset :  std_logic;
	SIGNAL ready :  std_logic;

BEGIN

	uut: ARS_rsacypher PORT MAP(
		indata => indata,
		inexp => inexp,
		inmod => inmod,
		cypher => cypher,
		clk => clk,
		ds => ds,
		reset => reset,
		ready => ready
	);


-- *** Test Bench - User Defined Section ***
	TB: PROCESS
	BEGIN
		wait for 120ns;
		reset <= '1';
		ds <= '0';
		wait for 20ns;
		wait until clk = '0';
		reset <= '0';
		wait until clk = '1';
		wait until clk = '0';
		--inexp <= x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001";
		--inexp <= 21789340966119291045314432534641202532740266679494864642379742093962117612319809219669273931607607861214081241256227427914086001225379063468332819468308212356077751884076761302314054656055360312570221352841005147503592134286229246963725459094556457331421004526308877633477209952149191344052218685160204715105191355183170454795905747626279346636011395174946384032654167498490215416634286862397602414656424535591397605573888224962313399362828588627807345215061836004345040558429385949651240843096176521766313185444868131902257530785588155477930469359255481573145685607784056994449421511113662704784792558507354925060519;
		inexp <=  x"192b7863caf59b10abd981c9ace9b88d3d3303d4ff7f3dfaf1d9f2e66090e7a91a0c621f6d88f0f20dbb8a3e60cdd644cfdb824553e46c005eb187ed3551c48ab90c6583421d5c9f90ce27ff9b76f3848dd866ee4ba4ce15167fbd3feda4cdced4230ee77736c3684aedf22e311594b2c409d0a183b0d0f99837bfe6fe9ede01";
		--inmod <=  23064945257292281727870978339468934825922468561893177588377650321255690350195208067466955625185006629763590496211713651839947130032069911035390515513973082829360541488534286899047787919981895536027493106058663141826265321575890316655519410552188910758981405732133455379422064526952626082517852182049524195378118440967128563456920250580707730892464377454506876576034962169619324118195349122945476969181614024480623086508459244181159254587208137962499274656454733972242297911580875021750217468245962574382071784183383565101930165596565611843030035142189452140462641597579988382551118268259060426206137653643644583749163;
		inmod <=  x"cc2d8d552f9b4c98b287dcdd63621e324fab5d61dc3381b38084fb9b1764ddfffda38ae0e7744670b36640e47f431d95a981210344d91dd7b74e8231a955c5c81a765dfb33c0312056a5c2a70e84a9f39f4e7297eee5e56158c8d14e0168047ea3f19d8971cc4818b3805d546f2163cab6916273db6f3a3ba005750e36b71151";
		indata <= x"1234567800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000087654321"; 
		--indata<= x"0011223300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000332211"; 
		--indata<=  x"9eeba2dedc2bd0ffefe0e51cc1e84e263c4b25f12328b9486fbd50ab1f5a8e4e74ad556f3a06f4a722cc01cc92e6aac7f7bad4ee19a496832f7027ca822b73625a572b16fcb5fe393347fef603bdf3eaa79b46bb833a5f4c393c6ddc612c2504b896a7b075ec821e79d7bf1d4d3c9cfca41c416f978c50be9188c156ae3af4e2";
		wait until clk = '1';
		wait for 2ns;
		ds <= '1';
		wait until ready = '0';
		ds <= '0';
		wait until ready = '1';
		wait;
		--$display("The encrypted data is :%h", cypher);
-- decrypt exponent		inexp <= x"02d80e39";
	END PROCESS;


   ClkGen : PROCESS
   BEGIN
      wait for 5300ps; -- will wait forever
		if clk = '1' then
			clk <= '0';
		else
			clk <= '1';
		end if;
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
